
`timescale 1ns / 1ps

module tb_N7_array_multiplier;

    // Parameters
    
    parameter N = 7;
    
     
    // Inputs
    
    reg  [6:0] A;
    
    reg  [6:0] B;
    
    
    // Outputs
    
    wire   P;
    
    
    // Instantiate the Unit Under Test (UUT)
    array_multiplier  #( N ) uut (
        
        .A(A),
        
        .B(B),
        
        
        .P(P)
        
    );

    // Clock generation 
    

    
    
    initial begin
        // Initialize Inputs
        
        A = 0;
        
        B = 0;
        
    
        // Wait for global reset
        #100;
    
        // Stimuli
        
        #10 A = 7'b1100001; B = 7'b0011000; // Expected: {'P': 2328}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100001; B = 7'b0011000; | Outputs: P=%b | Expected: P=%d",
                 0,
                 
                 P
                 , 
                 
                 2328
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100000; B = 7'b1110010; // Expected: {'P': 3648}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100000; B = 7'b1110010; | Outputs: P=%b | Expected: P=%d",
                 1,
                 
                 P
                 , 
                 
                 3648
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100011; B = 7'b1001111; // Expected: {'P': 7821}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100011; B = 7'b1001111; | Outputs: P=%b | Expected: P=%d",
                 2,
                 
                 P
                 , 
                 
                 7821
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110001; B = 7'b0110101; // Expected: {'P': 5989}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110001; B = 7'b0110101; | Outputs: P=%b | Expected: P=%d",
                 3,
                 
                 P
                 , 
                 
                 5989
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000011; B = 7'b1010011; // Expected: {'P': 249}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000011; B = 7'b1010011; | Outputs: P=%b | Expected: P=%d",
                 4,
                 
                 P
                 , 
                 
                 249
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101111; B = 7'b1000100; // Expected: {'P': 7548}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101111; B = 7'b1000100; | Outputs: P=%b | Expected: P=%d",
                 5,
                 
                 P
                 , 
                 
                 7548
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100010; B = 7'b1110100; // Expected: {'P': 3944}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100010; B = 7'b1110100; | Outputs: P=%b | Expected: P=%d",
                 6,
                 
                 P
                 , 
                 
                 3944
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001001; B = 7'b0100001; // Expected: {'P': 297}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001001; B = 7'b0100001; | Outputs: P=%b | Expected: P=%d",
                 7,
                 
                 P
                 , 
                 
                 297
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110101; B = 7'b1111110; // Expected: {'P': 6678}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110101; B = 7'b1111110; | Outputs: P=%b | Expected: P=%d",
                 8,
                 
                 P
                 , 
                 
                 6678
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011100; B = 7'b0001111; // Expected: {'P': 420}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011100; B = 7'b0001111; | Outputs: P=%b | Expected: P=%d",
                 9,
                 
                 P
                 , 
                 
                 420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100001; B = 7'b1010001; // Expected: {'P': 2673}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100001; B = 7'b1010001; | Outputs: P=%b | Expected: P=%d",
                 10,
                 
                 P
                 , 
                 
                 2673
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111111; B = 7'b0010111; // Expected: {'P': 2921}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111111; B = 7'b0010111; | Outputs: P=%b | Expected: P=%d",
                 11,
                 
                 P
                 , 
                 
                 2921
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000011; B = 7'b1011101; // Expected: {'P': 6231}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000011; B = 7'b1011101; | Outputs: P=%b | Expected: P=%d",
                 12,
                 
                 P
                 , 
                 
                 6231
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010100; B = 7'b0100001; // Expected: {'P': 660}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010100; B = 7'b0100001; | Outputs: P=%b | Expected: P=%d",
                 13,
                 
                 P
                 , 
                 
                 660
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010101; B = 7'b1011111; // Expected: {'P': 8075}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010101; B = 7'b1011111; | Outputs: P=%b | Expected: P=%d",
                 14,
                 
                 P
                 , 
                 
                 8075
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111000; B = 7'b1100010; // Expected: {'P': 5488}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111000; B = 7'b1100010; | Outputs: P=%b | Expected: P=%d",
                 15,
                 
                 P
                 , 
                 
                 5488
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000110; B = 7'b0111011; // Expected: {'P': 354}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000110; B = 7'b0111011; | Outputs: P=%b | Expected: P=%d",
                 16,
                 
                 P
                 , 
                 
                 354
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111101; B = 7'b1011011; // Expected: {'P': 5551}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111101; B = 7'b1011011; | Outputs: P=%b | Expected: P=%d",
                 17,
                 
                 P
                 , 
                 
                 5551
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011000; B = 7'b1110111; // Expected: {'P': 2856}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011000; B = 7'b1110111; | Outputs: P=%b | Expected: P=%d",
                 18,
                 
                 P
                 , 
                 
                 2856
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110011; B = 7'b0110111; // Expected: {'P': 6325}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110011; B = 7'b0110111; | Outputs: P=%b | Expected: P=%d",
                 19,
                 
                 P
                 , 
                 
                 6325
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111110; B = 7'b1011001; // Expected: {'P': 5518}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111110; B = 7'b1011001; | Outputs: P=%b | Expected: P=%d",
                 20,
                 
                 P
                 , 
                 
                 5518
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100000; B = 7'b0001111; // Expected: {'P': 1440}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100000; B = 7'b0001111; | Outputs: P=%b | Expected: P=%d",
                 21,
                 
                 P
                 , 
                 
                 1440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000011; B = 7'b0000110; // Expected: {'P': 402}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000011; B = 7'b0000110; | Outputs: P=%b | Expected: P=%d",
                 22,
                 
                 P
                 , 
                 
                 402
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011000; B = 7'b0110011; // Expected: {'P': 1224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011000; B = 7'b0110011; | Outputs: P=%b | Expected: P=%d",
                 23,
                 
                 P
                 , 
                 
                 1224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010000; B = 7'b0011111; // Expected: {'P': 496}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010000; B = 7'b0011111; | Outputs: P=%b | Expected: P=%d",
                 24,
                 
                 P
                 , 
                 
                 496
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011110; B = 7'b1001101; // Expected: {'P': 7238}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011110; B = 7'b1001101; | Outputs: P=%b | Expected: P=%d",
                 25,
                 
                 P
                 , 
                 
                 7238
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011101; B = 7'b0001001; // Expected: {'P': 261}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011101; B = 7'b0001001; | Outputs: P=%b | Expected: P=%d",
                 26,
                 
                 P
                 , 
                 
                 261
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110101; B = 7'b0101101; // Expected: {'P': 2385}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110101; B = 7'b0101101; | Outputs: P=%b | Expected: P=%d",
                 27,
                 
                 P
                 , 
                 
                 2385
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111100; B = 7'b1100110; // Expected: {'P': 6120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111100; B = 7'b1100110; | Outputs: P=%b | Expected: P=%d",
                 28,
                 
                 P
                 , 
                 
                 6120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001011; B = 7'b0000110; // Expected: {'P': 66}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001011; B = 7'b0000110; | Outputs: P=%b | Expected: P=%d",
                 29,
                 
                 P
                 , 
                 
                 66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011000; B = 7'b0011110; // Expected: {'P': 720}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011000; B = 7'b0011110; | Outputs: P=%b | Expected: P=%d",
                 30,
                 
                 P
                 , 
                 
                 720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111011; B = 7'b1001110; // Expected: {'P': 9594}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111011; B = 7'b1001110; | Outputs: P=%b | Expected: P=%d",
                 31,
                 
                 P
                 , 
                 
                 9594
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100000; B = 7'b1100101; // Expected: {'P': 3232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100000; B = 7'b1100101; | Outputs: P=%b | Expected: P=%d",
                 32,
                 
                 P
                 , 
                 
                 3232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010010; B = 7'b1101111; // Expected: {'P': 9102}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010010; B = 7'b1101111; | Outputs: P=%b | Expected: P=%d",
                 33,
                 
                 P
                 , 
                 
                 9102
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000010; B = 7'b0011111; // Expected: {'P': 2046}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000010; B = 7'b0011111; | Outputs: P=%b | Expected: P=%d",
                 34,
                 
                 P
                 , 
                 
                 2046
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000110; B = 7'b1010011; // Expected: {'P': 498}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000110; B = 7'b1010011; | Outputs: P=%b | Expected: P=%d",
                 35,
                 
                 P
                 , 
                 
                 498
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100011; B = 7'b0001100; // Expected: {'P': 1188}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100011; B = 7'b0001100; | Outputs: P=%b | Expected: P=%d",
                 36,
                 
                 P
                 , 
                 
                 1188
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100010; B = 7'b0010100; // Expected: {'P': 1960}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100010; B = 7'b0010100; | Outputs: P=%b | Expected: P=%d",
                 37,
                 
                 P
                 , 
                 
                 1960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110101; B = 7'b0001011; // Expected: {'P': 1287}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110101; B = 7'b0001011; | Outputs: P=%b | Expected: P=%d",
                 38,
                 
                 P
                 , 
                 
                 1287
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110100; B = 7'b0011001; // Expected: {'P': 2900}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110100; B = 7'b0011001; | Outputs: P=%b | Expected: P=%d",
                 39,
                 
                 P
                 , 
                 
                 2900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110000; B = 7'b1101100; // Expected: {'P': 5184}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110000; B = 7'b1101100; | Outputs: P=%b | Expected: P=%d",
                 40,
                 
                 P
                 , 
                 
                 5184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110001; B = 7'b1001100; // Expected: {'P': 8588}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110001; B = 7'b1001100; | Outputs: P=%b | Expected: P=%d",
                 41,
                 
                 P
                 , 
                 
                 8588
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000110; B = 7'b1101111; // Expected: {'P': 666}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000110; B = 7'b1101111; | Outputs: P=%b | Expected: P=%d",
                 42,
                 
                 P
                 , 
                 
                 666
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110010; B = 7'b1010111; // Expected: {'P': 4350}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110010; B = 7'b1010111; | Outputs: P=%b | Expected: P=%d",
                 43,
                 
                 P
                 , 
                 
                 4350
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100111; B = 7'b1011010; // Expected: {'P': 9270}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100111; B = 7'b1011010; | Outputs: P=%b | Expected: P=%d",
                 44,
                 
                 P
                 , 
                 
                 9270
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000011; B = 7'b1011001; // Expected: {'P': 5963}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000011; B = 7'b1011001; | Outputs: P=%b | Expected: P=%d",
                 45,
                 
                 P
                 , 
                 
                 5963
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101100; B = 7'b0110011; // Expected: {'P': 2244}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101100; B = 7'b0110011; | Outputs: P=%b | Expected: P=%d",
                 46,
                 
                 P
                 , 
                 
                 2244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000100; B = 7'b1101000; // Expected: {'P': 416}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000100; B = 7'b1101000; | Outputs: P=%b | Expected: P=%d",
                 47,
                 
                 P
                 , 
                 
                 416
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010101; B = 7'b1000101; // Expected: {'P': 1449}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010101; B = 7'b1000101; | Outputs: P=%b | Expected: P=%d",
                 48,
                 
                 P
                 , 
                 
                 1449
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100101; B = 7'b1000100; // Expected: {'P': 6868}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100101; B = 7'b1000100; | Outputs: P=%b | Expected: P=%d",
                 49,
                 
                 P
                 , 
                 
                 6868
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101101; B = 7'b0010100; // Expected: {'P': 2180}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101101; B = 7'b0010100; | Outputs: P=%b | Expected: P=%d",
                 50,
                 
                 P
                 , 
                 
                 2180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110010; B = 7'b1011001; // Expected: {'P': 10146}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110010; B = 7'b1011001; | Outputs: P=%b | Expected: P=%d",
                 51,
                 
                 P
                 , 
                 
                 10146
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011011; B = 7'b1100111; // Expected: {'P': 9373}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011011; B = 7'b1100111; | Outputs: P=%b | Expected: P=%d",
                 52,
                 
                 P
                 , 
                 
                 9373
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010001; B = 7'b1111011; // Expected: {'P': 2091}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010001; B = 7'b1111011; | Outputs: P=%b | Expected: P=%d",
                 53,
                 
                 P
                 , 
                 
                 2091
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010110; B = 7'b0000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010110; B = 7'b0000000; | Outputs: P=%b | Expected: P=%d",
                 54,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001011; B = 7'b0000001; // Expected: {'P': 11}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001011; B = 7'b0000001; | Outputs: P=%b | Expected: P=%d",
                 55,
                 
                 P
                 , 
                 
                 11
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000011; B = 7'b1111100; // Expected: {'P': 8308}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000011; B = 7'b1111100; | Outputs: P=%b | Expected: P=%d",
                 56,
                 
                 P
                 , 
                 
                 8308
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001110; B = 7'b0111011; // Expected: {'P': 826}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001110; B = 7'b0111011; | Outputs: P=%b | Expected: P=%d",
                 57,
                 
                 P
                 , 
                 
                 826
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101000; B = 7'b1010011; // Expected: {'P': 8632}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101000; B = 7'b1010011; | Outputs: P=%b | Expected: P=%d",
                 58,
                 
                 P
                 , 
                 
                 8632
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011001; B = 7'b1101111; // Expected: {'P': 2775}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011001; B = 7'b1101111; | Outputs: P=%b | Expected: P=%d",
                 59,
                 
                 P
                 , 
                 
                 2775
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001111; B = 7'b0001110; // Expected: {'P': 1106}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001111; B = 7'b0001110; | Outputs: P=%b | Expected: P=%d",
                 60,
                 
                 P
                 , 
                 
                 1106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100111; B = 7'b1101001; // Expected: {'P': 10815}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100111; B = 7'b1101001; | Outputs: P=%b | Expected: P=%d",
                 61,
                 
                 P
                 , 
                 
                 10815
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010110; B = 7'b0101000; // Expected: {'P': 880}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010110; B = 7'b0101000; | Outputs: P=%b | Expected: P=%d",
                 62,
                 
                 P
                 , 
                 
                 880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110110; B = 7'b1010110; // Expected: {'P': 4644}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110110; B = 7'b1010110; | Outputs: P=%b | Expected: P=%d",
                 63,
                 
                 P
                 , 
                 
                 4644
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100000; B = 7'b0111100; // Expected: {'P': 1920}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100000; B = 7'b0111100; | Outputs: P=%b | Expected: P=%d",
                 64,
                 
                 P
                 , 
                 
                 1920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010101; B = 7'b0100010; // Expected: {'P': 714}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010101; B = 7'b0100010; | Outputs: P=%b | Expected: P=%d",
                 65,
                 
                 P
                 , 
                 
                 714
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000011; B = 7'b1011010; // Expected: {'P': 6030}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000011; B = 7'b1011010; | Outputs: P=%b | Expected: P=%d",
                 66,
                 
                 P
                 , 
                 
                 6030
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100111; B = 7'b0111101; // Expected: {'P': 6283}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100111; B = 7'b0111101; | Outputs: P=%b | Expected: P=%d",
                 67,
                 
                 P
                 , 
                 
                 6283
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000110; B = 7'b0011111; // Expected: {'P': 2170}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000110; B = 7'b0011111; | Outputs: P=%b | Expected: P=%d",
                 68,
                 
                 P
                 , 
                 
                 2170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111110; B = 7'b1101100; // Expected: {'P': 13608}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111110; B = 7'b1101100; | Outputs: P=%b | Expected: P=%d",
                 69,
                 
                 P
                 , 
                 
                 13608
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001001; B = 7'b0001011; // Expected: {'P': 803}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001001; B = 7'b0001011; | Outputs: P=%b | Expected: P=%d",
                 70,
                 
                 P
                 , 
                 
                 803
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001011; B = 7'b1111111; // Expected: {'P': 1397}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001011; B = 7'b1111111; | Outputs: P=%b | Expected: P=%d",
                 71,
                 
                 P
                 , 
                 
                 1397
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001011; B = 7'b0100101; // Expected: {'P': 407}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001011; B = 7'b0100101; | Outputs: P=%b | Expected: P=%d",
                 72,
                 
                 P
                 , 
                 
                 407
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000000; B = 7'b1001000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000000; B = 7'b1001000; | Outputs: P=%b | Expected: P=%d",
                 73,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101110; B = 7'b1100110; // Expected: {'P': 11220}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101110; B = 7'b1100110; | Outputs: P=%b | Expected: P=%d",
                 74,
                 
                 P
                 , 
                 
                 11220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011110; B = 7'b0011101; // Expected: {'P': 870}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011110; B = 7'b0011101; | Outputs: P=%b | Expected: P=%d",
                 75,
                 
                 P
                 , 
                 
                 870
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010001; B = 7'b1110010; // Expected: {'P': 9234}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010001; B = 7'b1110010; | Outputs: P=%b | Expected: P=%d",
                 76,
                 
                 P
                 , 
                 
                 9234
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010110; B = 7'b0111101; // Expected: {'P': 1342}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010110; B = 7'b0111101; | Outputs: P=%b | Expected: P=%d",
                 77,
                 
                 P
                 , 
                 
                 1342
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101000; B = 7'b0100001; // Expected: {'P': 3432}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101000; B = 7'b0100001; | Outputs: P=%b | Expected: P=%d",
                 78,
                 
                 P
                 , 
                 
                 3432
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111001; B = 7'b0010111; // Expected: {'P': 1311}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111001; B = 7'b0010111; | Outputs: P=%b | Expected: P=%d",
                 79,
                 
                 P
                 , 
                 
                 1311
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100110; B = 7'b1111000; // Expected: {'P': 12240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100110; B = 7'b1111000; | Outputs: P=%b | Expected: P=%d",
                 80,
                 
                 P
                 , 
                 
                 12240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110001; B = 7'b0001011; // Expected: {'P': 1243}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110001; B = 7'b0001011; | Outputs: P=%b | Expected: P=%d",
                 81,
                 
                 P
                 , 
                 
                 1243
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011100; B = 7'b1101100; // Expected: {'P': 3024}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011100; B = 7'b1101100; | Outputs: P=%b | Expected: P=%d",
                 82,
                 
                 P
                 , 
                 
                 3024
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010100; B = 7'b0101001; // Expected: {'P': 3444}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010100; B = 7'b0101001; | Outputs: P=%b | Expected: P=%d",
                 83,
                 
                 P
                 , 
                 
                 3444
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100001; B = 7'b0001011; // Expected: {'P': 363}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100001; B = 7'b0001011; | Outputs: P=%b | Expected: P=%d",
                 84,
                 
                 P
                 , 
                 
                 363
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100100; B = 7'b0010001; // Expected: {'P': 1700}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100100; B = 7'b0010001; | Outputs: P=%b | Expected: P=%d",
                 85,
                 
                 P
                 , 
                 
                 1700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100001; B = 7'b1100101; // Expected: {'P': 9797}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100001; B = 7'b1100101; | Outputs: P=%b | Expected: P=%d",
                 86,
                 
                 P
                 , 
                 
                 9797
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000111; B = 7'b0010011; // Expected: {'P': 133}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000111; B = 7'b0010011; | Outputs: P=%b | Expected: P=%d",
                 87,
                 
                 P
                 , 
                 
                 133
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011011; B = 7'b0001101; // Expected: {'P': 351}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011011; B = 7'b0001101; | Outputs: P=%b | Expected: P=%d",
                 88,
                 
                 P
                 , 
                 
                 351
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100100; B = 7'b0000100; // Expected: {'P': 144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100100; B = 7'b0000100; | Outputs: P=%b | Expected: P=%d",
                 89,
                 
                 P
                 , 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000101; B = 7'b1011001; // Expected: {'P': 445}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000101; B = 7'b1011001; | Outputs: P=%b | Expected: P=%d",
                 90,
                 
                 P
                 , 
                 
                 445
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011010; B = 7'b1011110; // Expected: {'P': 2444}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011010; B = 7'b1011110; | Outputs: P=%b | Expected: P=%d",
                 91,
                 
                 P
                 , 
                 
                 2444
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110001; B = 7'b0010000; // Expected: {'P': 1808}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110001; B = 7'b0010000; | Outputs: P=%b | Expected: P=%d",
                 92,
                 
                 P
                 , 
                 
                 1808
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000001; B = 7'b1000111; // Expected: {'P': 71}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000001; B = 7'b1000111; | Outputs: P=%b | Expected: P=%d",
                 93,
                 
                 P
                 , 
                 
                 71
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000001; B = 7'b0100011; // Expected: {'P': 2275}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000001; B = 7'b0100011; | Outputs: P=%b | Expected: P=%d",
                 94,
                 
                 P
                 , 
                 
                 2275
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000011; B = 7'b0001010; // Expected: {'P': 670}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000011; B = 7'b0001010; | Outputs: P=%b | Expected: P=%d",
                 95,
                 
                 P
                 , 
                 
                 670
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110100; B = 7'b0011111; // Expected: {'P': 1612}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110100; B = 7'b0011111; | Outputs: P=%b | Expected: P=%d",
                 96,
                 
                 P
                 , 
                 
                 1612
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000111; B = 7'b1001011; // Expected: {'P': 525}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000111; B = 7'b1001011; | Outputs: P=%b | Expected: P=%d",
                 97,
                 
                 P
                 , 
                 
                 525
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011111; B = 7'b1110010; // Expected: {'P': 3534}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011111; B = 7'b1110010; | Outputs: P=%b | Expected: P=%d",
                 98,
                 
                 P
                 , 
                 
                 3534
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110110; B = 7'b0000010; // Expected: {'P': 236}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110110; B = 7'b0000010; | Outputs: P=%b | Expected: P=%d",
                 99,
                 
                 P
                 , 
                 
                 236
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111101; B = 7'b1110111; // Expected: {'P': 7259}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111101; B = 7'b1110111; | Outputs: P=%b | Expected: P=%d",
                 100,
                 
                 P
                 , 
                 
                 7259
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111101; B = 7'b0111111; // Expected: {'P': 7875}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111101; B = 7'b0111111; | Outputs: P=%b | Expected: P=%d",
                 101,
                 
                 P
                 , 
                 
                 7875
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001100; B = 7'b0101001; // Expected: {'P': 492}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001100; B = 7'b0101001; | Outputs: P=%b | Expected: P=%d",
                 102,
                 
                 P
                 , 
                 
                 492
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011011; B = 7'b0000100; // Expected: {'P': 108}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011011; B = 7'b0000100; | Outputs: P=%b | Expected: P=%d",
                 103,
                 
                 P
                 , 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010110; B = 7'b0001110; // Expected: {'P': 1204}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010110; B = 7'b0001110; | Outputs: P=%b | Expected: P=%d",
                 104,
                 
                 P
                 , 
                 
                 1204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000100; B = 7'b1100100; // Expected: {'P': 6800}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000100; B = 7'b1100100; | Outputs: P=%b | Expected: P=%d",
                 105,
                 
                 P
                 , 
                 
                 6800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011111; B = 7'b0010101; // Expected: {'P': 651}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011111; B = 7'b0010101; | Outputs: P=%b | Expected: P=%d",
                 106,
                 
                 P
                 , 
                 
                 651
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010000; B = 7'b1101100; // Expected: {'P': 1728}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010000; B = 7'b1101100; | Outputs: P=%b | Expected: P=%d",
                 107,
                 
                 P
                 , 
                 
                 1728
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110110; B = 7'b1001110; // Expected: {'P': 9204}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110110; B = 7'b1001110; | Outputs: P=%b | Expected: P=%d",
                 108,
                 
                 P
                 , 
                 
                 9204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010001; B = 7'b1110111; // Expected: {'P': 2023}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010001; B = 7'b1110111; | Outputs: P=%b | Expected: P=%d",
                 109,
                 
                 P
                 , 
                 
                 2023
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101010; B = 7'b1010000; // Expected: {'P': 8480}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101010; B = 7'b1010000; | Outputs: P=%b | Expected: P=%d",
                 110,
                 
                 P
                 , 
                 
                 8480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101000; B = 7'b1110101; // Expected: {'P': 12168}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101000; B = 7'b1110101; | Outputs: P=%b | Expected: P=%d",
                 111,
                 
                 P
                 , 
                 
                 12168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010100; B = 7'b0100100; // Expected: {'P': 720}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010100; B = 7'b0100100; | Outputs: P=%b | Expected: P=%d",
                 112,
                 
                 P
                 , 
                 
                 720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001010; B = 7'b0000111; // Expected: {'P': 70}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001010; B = 7'b0000111; | Outputs: P=%b | Expected: P=%d",
                 113,
                 
                 P
                 , 
                 
                 70
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000100; B = 7'b0001111; // Expected: {'P': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000100; B = 7'b0001111; | Outputs: P=%b | Expected: P=%d",
                 114,
                 
                 P
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001011; B = 7'b0101001; // Expected: {'P': 451}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001011; B = 7'b0101001; | Outputs: P=%b | Expected: P=%d",
                 115,
                 
                 P
                 , 
                 
                 451
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111010; B = 7'b0111001; // Expected: {'P': 3306}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111010; B = 7'b0111001; | Outputs: P=%b | Expected: P=%d",
                 116,
                 
                 P
                 , 
                 
                 3306
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010001; B = 7'b1111001; // Expected: {'P': 9801}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010001; B = 7'b1111001; | Outputs: P=%b | Expected: P=%d",
                 117,
                 
                 P
                 , 
                 
                 9801
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001101; B = 7'b0001001; // Expected: {'P': 693}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001101; B = 7'b0001001; | Outputs: P=%b | Expected: P=%d",
                 118,
                 
                 P
                 , 
                 
                 693
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101011; B = 7'b0100010; // Expected: {'P': 3638}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101011; B = 7'b0100010; | Outputs: P=%b | Expected: P=%d",
                 119,
                 
                 P
                 , 
                 
                 3638
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110001; B = 7'b1100110; // Expected: {'P': 11526}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110001; B = 7'b1100110; | Outputs: P=%b | Expected: P=%d",
                 120,
                 
                 P
                 , 
                 
                 11526
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010100; B = 7'b1100001; // Expected: {'P': 8148}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010100; B = 7'b1100001; | Outputs: P=%b | Expected: P=%d",
                 121,
                 
                 P
                 , 
                 
                 8148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010001; B = 7'b0011101; // Expected: {'P': 493}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010001; B = 7'b0011101; | Outputs: P=%b | Expected: P=%d",
                 122,
                 
                 P
                 , 
                 
                 493
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010111; B = 7'b0110100; // Expected: {'P': 1196}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010111; B = 7'b0110100; | Outputs: P=%b | Expected: P=%d",
                 123,
                 
                 P
                 , 
                 
                 1196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111100; B = 7'b0000100; // Expected: {'P': 496}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111100; B = 7'b0000100; | Outputs: P=%b | Expected: P=%d",
                 124,
                 
                 P
                 , 
                 
                 496
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111000; B = 7'b1000101; // Expected: {'P': 3864}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111000; B = 7'b1000101; | Outputs: P=%b | Expected: P=%d",
                 125,
                 
                 P
                 , 
                 
                 3864
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010000; B = 7'b1110010; // Expected: {'P': 1824}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010000; B = 7'b1110010; | Outputs: P=%b | Expected: P=%d",
                 126,
                 
                 P
                 , 
                 
                 1824
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011000; B = 7'b1001011; // Expected: {'P': 1800}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011000; B = 7'b1001011; | Outputs: P=%b | Expected: P=%d",
                 127,
                 
                 P
                 , 
                 
                 1800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011110; B = 7'b1011001; // Expected: {'P': 8366}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011110; B = 7'b1011001; | Outputs: P=%b | Expected: P=%d",
                 128,
                 
                 P
                 , 
                 
                 8366
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000111; B = 7'b0110001; // Expected: {'P': 343}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000111; B = 7'b0110001; | Outputs: P=%b | Expected: P=%d",
                 129,
                 
                 P
                 , 
                 
                 343
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001011; B = 7'b1010001; // Expected: {'P': 891}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001011; B = 7'b1010001; | Outputs: P=%b | Expected: P=%d",
                 130,
                 
                 P
                 , 
                 
                 891
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111111; B = 7'b1101001; // Expected: {'P': 13335}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111111; B = 7'b1101001; | Outputs: P=%b | Expected: P=%d",
                 131,
                 
                 P
                 , 
                 
                 13335
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001101; B = 7'b0010011; // Expected: {'P': 247}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001101; B = 7'b0010011; | Outputs: P=%b | Expected: P=%d",
                 132,
                 
                 P
                 , 
                 
                 247
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011101; B = 7'b0010110; // Expected: {'P': 638}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011101; B = 7'b0010110; | Outputs: P=%b | Expected: P=%d",
                 133,
                 
                 P
                 , 
                 
                 638
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011010; B = 7'b1111001; // Expected: {'P': 3146}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011010; B = 7'b1111001; | Outputs: P=%b | Expected: P=%d",
                 134,
                 
                 P
                 , 
                 
                 3146
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001011; B = 7'b1111111; // Expected: {'P': 9525}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001011; B = 7'b1111111; | Outputs: P=%b | Expected: P=%d",
                 135,
                 
                 P
                 , 
                 
                 9525
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100001; B = 7'b0011101; // Expected: {'P': 957}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100001; B = 7'b0011101; | Outputs: P=%b | Expected: P=%d",
                 136,
                 
                 P
                 , 
                 
                 957
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100101; B = 7'b0011110; // Expected: {'P': 1110}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100101; B = 7'b0011110; | Outputs: P=%b | Expected: P=%d",
                 137,
                 
                 P
                 , 
                 
                 1110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101100; B = 7'b0110100; // Expected: {'P': 5616}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101100; B = 7'b0110100; | Outputs: P=%b | Expected: P=%d",
                 138,
                 
                 P
                 , 
                 
                 5616
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001010; B = 7'b0011110; // Expected: {'P': 2220}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001010; B = 7'b0011110; | Outputs: P=%b | Expected: P=%d",
                 139,
                 
                 P
                 , 
                 
                 2220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110010; B = 7'b1110001; // Expected: {'P': 5650}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110010; B = 7'b1110001; | Outputs: P=%b | Expected: P=%d",
                 140,
                 
                 P
                 , 
                 
                 5650
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011010; B = 7'b0110111; // Expected: {'P': 1430}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011010; B = 7'b0110111; | Outputs: P=%b | Expected: P=%d",
                 141,
                 
                 P
                 , 
                 
                 1430
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010011; B = 7'b1100011; // Expected: {'P': 1881}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010011; B = 7'b1100011; | Outputs: P=%b | Expected: P=%d",
                 142,
                 
                 P
                 , 
                 
                 1881
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101011; B = 7'b0100100; // Expected: {'P': 1548}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101011; B = 7'b0100100; | Outputs: P=%b | Expected: P=%d",
                 143,
                 
                 P
                 , 
                 
                 1548
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100100; B = 7'b1101010; // Expected: {'P': 10600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100100; B = 7'b1101010; | Outputs: P=%b | Expected: P=%d",
                 144,
                 
                 P
                 , 
                 
                 10600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100011; B = 7'b0110000; // Expected: {'P': 4752}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100011; B = 7'b0110000; | Outputs: P=%b | Expected: P=%d",
                 145,
                 
                 P
                 , 
                 
                 4752
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000101; B = 7'b0111001; // Expected: {'P': 285}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000101; B = 7'b0111001; | Outputs: P=%b | Expected: P=%d",
                 146,
                 
                 P
                 , 
                 
                 285
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001101; B = 7'b0001101; // Expected: {'P': 169}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001101; B = 7'b0001101; | Outputs: P=%b | Expected: P=%d",
                 147,
                 
                 P
                 , 
                 
                 169
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001110; B = 7'b0111011; // Expected: {'P': 4602}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001110; B = 7'b0111011; | Outputs: P=%b | Expected: P=%d",
                 148,
                 
                 P
                 , 
                 
                 4602
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110010; B = 7'b1100100; // Expected: {'P': 11400}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110010; B = 7'b1100100; | Outputs: P=%b | Expected: P=%d",
                 149,
                 
                 P
                 , 
                 
                 11400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101110; B = 7'b0011111; // Expected: {'P': 1426}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101110; B = 7'b0011111; | Outputs: P=%b | Expected: P=%d",
                 150,
                 
                 P
                 , 
                 
                 1426
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110101; B = 7'b0010001; // Expected: {'P': 901}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110101; B = 7'b0010001; | Outputs: P=%b | Expected: P=%d",
                 151,
                 
                 P
                 , 
                 
                 901
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010101; B = 7'b1100011; // Expected: {'P': 2079}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010101; B = 7'b1100011; | Outputs: P=%b | Expected: P=%d",
                 152,
                 
                 P
                 , 
                 
                 2079
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001101; B = 7'b1100010; // Expected: {'P': 7546}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001101; B = 7'b1100010; | Outputs: P=%b | Expected: P=%d",
                 153,
                 
                 P
                 , 
                 
                 7546
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110001; B = 7'b0110111; // Expected: {'P': 2695}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110001; B = 7'b0110111; | Outputs: P=%b | Expected: P=%d",
                 154,
                 
                 P
                 , 
                 
                 2695
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010101; B = 7'b0100001; // Expected: {'P': 693}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010101; B = 7'b0100001; | Outputs: P=%b | Expected: P=%d",
                 155,
                 
                 P
                 , 
                 
                 693
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010111; B = 7'b0000001; // Expected: {'P': 23}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010111; B = 7'b0000001; | Outputs: P=%b | Expected: P=%d",
                 156,
                 
                 P
                 , 
                 
                 23
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100101; B = 7'b0110000; // Expected: {'P': 4848}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100101; B = 7'b0110000; | Outputs: P=%b | Expected: P=%d",
                 157,
                 
                 P
                 , 
                 
                 4848
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100010; B = 7'b0100011; // Expected: {'P': 1190}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100010; B = 7'b0100011; | Outputs: P=%b | Expected: P=%d",
                 158,
                 
                 P
                 , 
                 
                 1190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001110; B = 7'b1110100; // Expected: {'P': 1624}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001110; B = 7'b1110100; | Outputs: P=%b | Expected: P=%d",
                 159,
                 
                 P
                 , 
                 
                 1624
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110100; B = 7'b1010100; // Expected: {'P': 4368}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110100; B = 7'b1010100; | Outputs: P=%b | Expected: P=%d",
                 160,
                 
                 P
                 , 
                 
                 4368
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110111; B = 7'b1011011; // Expected: {'P': 10829}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110111; B = 7'b1011011; | Outputs: P=%b | Expected: P=%d",
                 161,
                 
                 P
                 , 
                 
                 10829
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101111; B = 7'b0101000; // Expected: {'P': 1880}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101111; B = 7'b0101000; | Outputs: P=%b | Expected: P=%d",
                 162,
                 
                 P
                 , 
                 
                 1880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110101; B = 7'b0011000; // Expected: {'P': 2808}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110101; B = 7'b0011000; | Outputs: P=%b | Expected: P=%d",
                 163,
                 
                 P
                 , 
                 
                 2808
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000000; B = 7'b1111110; // Expected: {'P': 8064}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000000; B = 7'b1111110; | Outputs: P=%b | Expected: P=%d",
                 164,
                 
                 P
                 , 
                 
                 8064
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100001; B = 7'b0110111; // Expected: {'P': 1815}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100001; B = 7'b0110111; | Outputs: P=%b | Expected: P=%d",
                 165,
                 
                 P
                 , 
                 
                 1815
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001011; B = 7'b1101000; // Expected: {'P': 1144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001011; B = 7'b1101000; | Outputs: P=%b | Expected: P=%d",
                 166,
                 
                 P
                 , 
                 
                 1144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110001; B = 7'b0011111; // Expected: {'P': 3503}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110001; B = 7'b0011111; | Outputs: P=%b | Expected: P=%d",
                 167,
                 
                 P
                 , 
                 
                 3503
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101001; B = 7'b0010100; // Expected: {'P': 2100}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101001; B = 7'b0010100; | Outputs: P=%b | Expected: P=%d",
                 168,
                 
                 P
                 , 
                 
                 2100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000011; B = 7'b1110101; // Expected: {'P': 7839}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000011; B = 7'b1110101; | Outputs: P=%b | Expected: P=%d",
                 169,
                 
                 P
                 , 
                 
                 7839
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001111; B = 7'b0001011; // Expected: {'P': 869}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001111; B = 7'b0001011; | Outputs: P=%b | Expected: P=%d",
                 170,
                 
                 P
                 , 
                 
                 869
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001010; B = 7'b1010110; // Expected: {'P': 6364}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001010; B = 7'b1010110; | Outputs: P=%b | Expected: P=%d",
                 171,
                 
                 P
                 , 
                 
                 6364
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111011; B = 7'b1100101; // Expected: {'P': 12423}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111011; B = 7'b1100101; | Outputs: P=%b | Expected: P=%d",
                 172,
                 
                 P
                 , 
                 
                 12423
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111010; B = 7'b0000101; // Expected: {'P': 290}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111010; B = 7'b0000101; | Outputs: P=%b | Expected: P=%d",
                 173,
                 
                 P
                 , 
                 
                 290
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011110; B = 7'b0000101; // Expected: {'P': 150}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011110; B = 7'b0000101; | Outputs: P=%b | Expected: P=%d",
                 174,
                 
                 P
                 , 
                 
                 150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100110; B = 7'b0101100; // Expected: {'P': 1672}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100110; B = 7'b0101100; | Outputs: P=%b | Expected: P=%d",
                 175,
                 
                 P
                 , 
                 
                 1672
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101101; B = 7'b1000000; // Expected: {'P': 6976}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101101; B = 7'b1000000; | Outputs: P=%b | Expected: P=%d",
                 176,
                 
                 P
                 , 
                 
                 6976
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110110; B = 7'b1101101; // Expected: {'P': 5886}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110110; B = 7'b1101101; | Outputs: P=%b | Expected: P=%d",
                 177,
                 
                 P
                 , 
                 
                 5886
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110111; B = 7'b1110011; // Expected: {'P': 13685}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110111; B = 7'b1110011; | Outputs: P=%b | Expected: P=%d",
                 178,
                 
                 P
                 , 
                 
                 13685
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001010; B = 7'b1111010; // Expected: {'P': 1220}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001010; B = 7'b1111010; | Outputs: P=%b | Expected: P=%d",
                 179,
                 
                 P
                 , 
                 
                 1220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100011; B = 7'b0111001; // Expected: {'P': 5643}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100011; B = 7'b0111001; | Outputs: P=%b | Expected: P=%d",
                 180,
                 
                 P
                 , 
                 
                 5643
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100010; B = 7'b1100101; // Expected: {'P': 3434}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100010; B = 7'b1100101; | Outputs: P=%b | Expected: P=%d",
                 181,
                 
                 P
                 , 
                 
                 3434
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010010; B = 7'b0010101; // Expected: {'P': 378}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010010; B = 7'b0010101; | Outputs: P=%b | Expected: P=%d",
                 182,
                 
                 P
                 , 
                 
                 378
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000111; B = 7'b1100000; // Expected: {'P': 672}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000111; B = 7'b1100000; | Outputs: P=%b | Expected: P=%d",
                 183,
                 
                 P
                 , 
                 
                 672
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011101; B = 7'b0000001; // Expected: {'P': 29}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011101; B = 7'b0000001; | Outputs: P=%b | Expected: P=%d",
                 184,
                 
                 P
                 , 
                 
                 29
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000101; B = 7'b1001101; // Expected: {'P': 5313}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000101; B = 7'b1001101; | Outputs: P=%b | Expected: P=%d",
                 185,
                 
                 P
                 , 
                 
                 5313
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010000; B = 7'b1100100; // Expected: {'P': 8000}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010000; B = 7'b1100100; | Outputs: P=%b | Expected: P=%d",
                 186,
                 
                 P
                 , 
                 
                 8000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101000; B = 7'b0010111; // Expected: {'P': 2392}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101000; B = 7'b0010111; | Outputs: P=%b | Expected: P=%d",
                 187,
                 
                 P
                 , 
                 
                 2392
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101010; B = 7'b1100010; // Expected: {'P': 4116}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101010; B = 7'b1100010; | Outputs: P=%b | Expected: P=%d",
                 188,
                 
                 P
                 , 
                 
                 4116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101100; B = 7'b1010001; // Expected: {'P': 8748}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101100; B = 7'b1010001; | Outputs: P=%b | Expected: P=%d",
                 189,
                 
                 P
                 , 
                 
                 8748
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001010; B = 7'b1000011; // Expected: {'P': 4958}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001010; B = 7'b1000011; | Outputs: P=%b | Expected: P=%d",
                 190,
                 
                 P
                 , 
                 
                 4958
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100010; B = 7'b1100001; // Expected: {'P': 3298}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100010; B = 7'b1100001; | Outputs: P=%b | Expected: P=%d",
                 191,
                 
                 P
                 , 
                 
                 3298
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101101; B = 7'b1011010; // Expected: {'P': 9810}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101101; B = 7'b1011010; | Outputs: P=%b | Expected: P=%d",
                 192,
                 
                 P
                 , 
                 
                 9810
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000101; B = 7'b0000011; // Expected: {'P': 15}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000101; B = 7'b0000011; | Outputs: P=%b | Expected: P=%d",
                 193,
                 
                 P
                 , 
                 
                 15
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001110; B = 7'b1101000; // Expected: {'P': 1456}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001110; B = 7'b1101000; | Outputs: P=%b | Expected: P=%d",
                 194,
                 
                 P
                 , 
                 
                 1456
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011010; B = 7'b0011010; // Expected: {'P': 2340}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011010; B = 7'b0011010; | Outputs: P=%b | Expected: P=%d",
                 195,
                 
                 P
                 , 
                 
                 2340
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110111; B = 7'b0001010; // Expected: {'P': 550}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110111; B = 7'b0001010; | Outputs: P=%b | Expected: P=%d",
                 196,
                 
                 P
                 , 
                 
                 550
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111110; B = 7'b0010011; // Expected: {'P': 2394}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111110; B = 7'b0010011; | Outputs: P=%b | Expected: P=%d",
                 197,
                 
                 P
                 , 
                 
                 2394
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101001; B = 7'b0111110; // Expected: {'P': 2542}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101001; B = 7'b0111110; | Outputs: P=%b | Expected: P=%d",
                 198,
                 
                 P
                 , 
                 
                 2542
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010001; B = 7'b1010000; // Expected: {'P': 6480}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010001; B = 7'b1010000; | Outputs: P=%b | Expected: P=%d",
                 199,
                 
                 P
                 , 
                 
                 6480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101011; B = 7'b1000010; // Expected: {'P': 2838}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101011; B = 7'b1000010; | Outputs: P=%b | Expected: P=%d",
                 200,
                 
                 P
                 , 
                 
                 2838
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001101; B = 7'b1110001; // Expected: {'P': 8701}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001101; B = 7'b1110001; | Outputs: P=%b | Expected: P=%d",
                 201,
                 
                 P
                 , 
                 
                 8701
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000001; B = 7'b1000110; // Expected: {'P': 4550}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000001; B = 7'b1000110; | Outputs: P=%b | Expected: P=%d",
                 202,
                 
                 P
                 , 
                 
                 4550
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000000; B = 7'b0010001; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000000; B = 7'b0010001; | Outputs: P=%b | Expected: P=%d",
                 203,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000001; B = 7'b1010101; // Expected: {'P': 85}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000001; B = 7'b1010101; | Outputs: P=%b | Expected: P=%d",
                 204,
                 
                 P
                 , 
                 
                 85
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010110; B = 7'b0100000; // Expected: {'P': 2752}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010110; B = 7'b0100000; | Outputs: P=%b | Expected: P=%d",
                 205,
                 
                 P
                 , 
                 
                 2752
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101111; B = 7'b1110000; // Expected: {'P': 5264}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101111; B = 7'b1110000; | Outputs: P=%b | Expected: P=%d",
                 206,
                 
                 P
                 , 
                 
                 5264
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101100; B = 7'b1010010; // Expected: {'P': 3608}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101100; B = 7'b1010010; | Outputs: P=%b | Expected: P=%d",
                 207,
                 
                 P
                 , 
                 
                 3608
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011101; B = 7'b1111100; // Expected: {'P': 11532}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011101; B = 7'b1111100; | Outputs: P=%b | Expected: P=%d",
                 208,
                 
                 P
                 , 
                 
                 11532
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011001; B = 7'b0010011; // Expected: {'P': 475}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011001; B = 7'b0010011; | Outputs: P=%b | Expected: P=%d",
                 209,
                 
                 P
                 , 
                 
                 475
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100011; B = 7'b1001101; // Expected: {'P': 2695}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100011; B = 7'b1001101; | Outputs: P=%b | Expected: P=%d",
                 210,
                 
                 P
                 , 
                 
                 2695
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110010; B = 7'b0000111; // Expected: {'P': 350}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110010; B = 7'b0000111; | Outputs: P=%b | Expected: P=%d",
                 211,
                 
                 P
                 , 
                 
                 350
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011000; B = 7'b1110010; // Expected: {'P': 10032}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011000; B = 7'b1110010; | Outputs: P=%b | Expected: P=%d",
                 212,
                 
                 P
                 , 
                 
                 10032
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010000; B = 7'b1010010; // Expected: {'P': 6560}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010000; B = 7'b1010010; | Outputs: P=%b | Expected: P=%d",
                 213,
                 
                 P
                 , 
                 
                 6560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101001; B = 7'b1000111; // Expected: {'P': 2911}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101001; B = 7'b1000111; | Outputs: P=%b | Expected: P=%d",
                 214,
                 
                 P
                 , 
                 
                 2911
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011101; B = 7'b0100010; // Expected: {'P': 986}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011101; B = 7'b0100010; | Outputs: P=%b | Expected: P=%d",
                 215,
                 
                 P
                 , 
                 
                 986
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110011; B = 7'b0100001; // Expected: {'P': 3795}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110011; B = 7'b0100001; | Outputs: P=%b | Expected: P=%d",
                 216,
                 
                 P
                 , 
                 
                 3795
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000010; B = 7'b1001001; // Expected: {'P': 146}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000010; B = 7'b1001001; | Outputs: P=%b | Expected: P=%d",
                 217,
                 
                 P
                 , 
                 
                 146
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101110; B = 7'b1000101; // Expected: {'P': 3174}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101110; B = 7'b1000101; | Outputs: P=%b | Expected: P=%d",
                 218,
                 
                 P
                 , 
                 
                 3174
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111111; B = 7'b1010001; // Expected: {'P': 10287}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111111; B = 7'b1010001; | Outputs: P=%b | Expected: P=%d",
                 219,
                 
                 P
                 , 
                 
                 10287
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011010; B = 7'b1010010; // Expected: {'P': 2132}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011010; B = 7'b1010010; | Outputs: P=%b | Expected: P=%d",
                 220,
                 
                 P
                 , 
                 
                 2132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001111; B = 7'b1001011; // Expected: {'P': 5925}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001111; B = 7'b1001011; | Outputs: P=%b | Expected: P=%d",
                 221,
                 
                 P
                 , 
                 
                 5925
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010100; B = 7'b1110011; // Expected: {'P': 9660}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010100; B = 7'b1110011; | Outputs: P=%b | Expected: P=%d",
                 222,
                 
                 P
                 , 
                 
                 9660
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110100; B = 7'b1101101; // Expected: {'P': 5668}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110100; B = 7'b1101101; | Outputs: P=%b | Expected: P=%d",
                 223,
                 
                 P
                 , 
                 
                 5668
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111001; B = 7'b1000011; // Expected: {'P': 8107}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111001; B = 7'b1000011; | Outputs: P=%b | Expected: P=%d",
                 224,
                 
                 P
                 , 
                 
                 8107
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110000; B = 7'b0010110; // Expected: {'P': 1056}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110000; B = 7'b0010110; | Outputs: P=%b | Expected: P=%d",
                 225,
                 
                 P
                 , 
                 
                 1056
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001111; B = 7'b1111000; // Expected: {'P': 9480}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001111; B = 7'b1111000; | Outputs: P=%b | Expected: P=%d",
                 226,
                 
                 P
                 , 
                 
                 9480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011000; B = 7'b0110000; // Expected: {'P': 1152}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011000; B = 7'b0110000; | Outputs: P=%b | Expected: P=%d",
                 227,
                 
                 P
                 , 
                 
                 1152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111000; B = 7'b0111001; // Expected: {'P': 6840}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111000; B = 7'b0111001; | Outputs: P=%b | Expected: P=%d",
                 228,
                 
                 P
                 , 
                 
                 6840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100010; B = 7'b0000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100010; B = 7'b0000000; | Outputs: P=%b | Expected: P=%d",
                 229,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000011; B = 7'b1010001; // Expected: {'P': 5427}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000011; B = 7'b1010001; | Outputs: P=%b | Expected: P=%d",
                 230,
                 
                 P
                 , 
                 
                 5427
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100000; B = 7'b1001010; // Expected: {'P': 2368}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100000; B = 7'b1001010; | Outputs: P=%b | Expected: P=%d",
                 231,
                 
                 P
                 , 
                 
                 2368
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111110; B = 7'b0101100; // Expected: {'P': 2728}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111110; B = 7'b0101100; | Outputs: P=%b | Expected: P=%d",
                 232,
                 
                 P
                 , 
                 
                 2728
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000101; B = 7'b0001101; // Expected: {'P': 897}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000101; B = 7'b0001101; | Outputs: P=%b | Expected: P=%d",
                 233,
                 
                 P
                 , 
                 
                 897
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101001; B = 7'b0000101; // Expected: {'P': 205}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101001; B = 7'b0000101; | Outputs: P=%b | Expected: P=%d",
                 234,
                 
                 P
                 , 
                 
                 205
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111001; B = 7'b1100110; // Expected: {'P': 5814}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111001; B = 7'b1100110; | Outputs: P=%b | Expected: P=%d",
                 235,
                 
                 P
                 , 
                 
                 5814
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010110; B = 7'b1001110; // Expected: {'P': 1716}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010110; B = 7'b1001110; | Outputs: P=%b | Expected: P=%d",
                 236,
                 
                 P
                 , 
                 
                 1716
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100111; B = 7'b1000101; // Expected: {'P': 7107}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100111; B = 7'b1000101; | Outputs: P=%b | Expected: P=%d",
                 237,
                 
                 P
                 , 
                 
                 7107
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101111; B = 7'b0000100; // Expected: {'P': 444}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101111; B = 7'b0000100; | Outputs: P=%b | Expected: P=%d",
                 238,
                 
                 P
                 , 
                 
                 444
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110100; B = 7'b1000000; // Expected: {'P': 3328}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110100; B = 7'b1000000; | Outputs: P=%b | Expected: P=%d",
                 239,
                 
                 P
                 , 
                 
                 3328
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101110; B = 7'b0000110; // Expected: {'P': 276}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101110; B = 7'b0000110; | Outputs: P=%b | Expected: P=%d",
                 240,
                 
                 P
                 , 
                 
                 276
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010111; B = 7'b1011100; // Expected: {'P': 2116}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010111; B = 7'b1011100; | Outputs: P=%b | Expected: P=%d",
                 241,
                 
                 P
                 , 
                 
                 2116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001101; B = 7'b0100100; // Expected: {'P': 2772}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001101; B = 7'b0100100; | Outputs: P=%b | Expected: P=%d",
                 242,
                 
                 P
                 , 
                 
                 2772
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001101; B = 7'b1110000; // Expected: {'P': 8624}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001101; B = 7'b1110000; | Outputs: P=%b | Expected: P=%d",
                 243,
                 
                 P
                 , 
                 
                 8624
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001111; B = 7'b1111011; // Expected: {'P': 9717}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001111; B = 7'b1111011; | Outputs: P=%b | Expected: P=%d",
                 244,
                 
                 P
                 , 
                 
                 9717
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111001; B = 7'b1001111; // Expected: {'P': 4503}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111001; B = 7'b1001111; | Outputs: P=%b | Expected: P=%d",
                 245,
                 
                 P
                 , 
                 
                 4503
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001011; B = 7'b0000010; // Expected: {'P': 22}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001011; B = 7'b0000010; | Outputs: P=%b | Expected: P=%d",
                 246,
                 
                 P
                 , 
                 
                 22
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011111; B = 7'b1000110; // Expected: {'P': 2170}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011111; B = 7'b1000110; | Outputs: P=%b | Expected: P=%d",
                 247,
                 
                 P
                 , 
                 
                 2170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110111; B = 7'b1001101; // Expected: {'P': 4235}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110111; B = 7'b1001101; | Outputs: P=%b | Expected: P=%d",
                 248,
                 
                 P
                 , 
                 
                 4235
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111010; B = 7'b1111000; // Expected: {'P': 14640}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111010; B = 7'b1111000; | Outputs: P=%b | Expected: P=%d",
                 249,
                 
                 P
                 , 
                 
                 14640
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001010; B = 7'b0101000; // Expected: {'P': 400}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001010; B = 7'b0101000; | Outputs: P=%b | Expected: P=%d",
                 250,
                 
                 P
                 , 
                 
                 400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010111; B = 7'b0110011; // Expected: {'P': 1173}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010111; B = 7'b0110011; | Outputs: P=%b | Expected: P=%d",
                 251,
                 
                 P
                 , 
                 
                 1173
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101111; B = 7'b1110110; // Expected: {'P': 13098}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101111; B = 7'b1110110; | Outputs: P=%b | Expected: P=%d",
                 252,
                 
                 P
                 , 
                 
                 13098
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001000; B = 7'b1001011; // Expected: {'P': 600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001000; B = 7'b1001011; | Outputs: P=%b | Expected: P=%d",
                 253,
                 
                 P
                 , 
                 
                 600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111000; B = 7'b1001111; // Expected: {'P': 9480}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111000; B = 7'b1001111; | Outputs: P=%b | Expected: P=%d",
                 254,
                 
                 P
                 , 
                 
                 9480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100101; B = 7'b1110000; // Expected: {'P': 4144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100101; B = 7'b1110000; | Outputs: P=%b | Expected: P=%d",
                 255,
                 
                 P
                 , 
                 
                 4144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111000; B = 7'b1100000; // Expected: {'P': 11520}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111000; B = 7'b1100000; | Outputs: P=%b | Expected: P=%d",
                 256,
                 
                 P
                 , 
                 
                 11520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101101; B = 7'b1101001; // Expected: {'P': 11445}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101101; B = 7'b1101001; | Outputs: P=%b | Expected: P=%d",
                 257,
                 
                 P
                 , 
                 
                 11445
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011111; B = 7'b0001011; // Expected: {'P': 341}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011111; B = 7'b0001011; | Outputs: P=%b | Expected: P=%d",
                 258,
                 
                 P
                 , 
                 
                 341
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100011; B = 7'b0010101; // Expected: {'P': 2079}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100011; B = 7'b0010101; | Outputs: P=%b | Expected: P=%d",
                 259,
                 
                 P
                 , 
                 
                 2079
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011101; B = 7'b1001011; // Expected: {'P': 6975}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011101; B = 7'b1001011; | Outputs: P=%b | Expected: P=%d",
                 260,
                 
                 P
                 , 
                 
                 6975
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000011; B = 7'b1101101; // Expected: {'P': 327}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000011; B = 7'b1101101; | Outputs: P=%b | Expected: P=%d",
                 261,
                 
                 P
                 , 
                 
                 327
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111111; B = 7'b0010000; // Expected: {'P': 1008}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111111; B = 7'b0010000; | Outputs: P=%b | Expected: P=%d",
                 262,
                 
                 P
                 , 
                 
                 1008
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010011; B = 7'b0100010; // Expected: {'P': 646}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010011; B = 7'b0100010; | Outputs: P=%b | Expected: P=%d",
                 263,
                 
                 P
                 , 
                 
                 646
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001011; B = 7'b1010101; // Expected: {'P': 935}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001011; B = 7'b1010101; | Outputs: P=%b | Expected: P=%d",
                 264,
                 
                 P
                 , 
                 
                 935
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101111; B = 7'b1110010; // Expected: {'P': 5358}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101111; B = 7'b1110010; | Outputs: P=%b | Expected: P=%d",
                 265,
                 
                 P
                 , 
                 
                 5358
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010001; B = 7'b1001001; // Expected: {'P': 1241}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010001; B = 7'b1001001; | Outputs: P=%b | Expected: P=%d",
                 266,
                 
                 P
                 , 
                 
                 1241
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000001; B = 7'b1011001; // Expected: {'P': 5785}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000001; B = 7'b1011001; | Outputs: P=%b | Expected: P=%d",
                 267,
                 
                 P
                 , 
                 
                 5785
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110111; B = 7'b1100001; // Expected: {'P': 11543}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110111; B = 7'b1100001; | Outputs: P=%b | Expected: P=%d",
                 268,
                 
                 P
                 , 
                 
                 11543
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101101; B = 7'b1011110; // Expected: {'P': 10246}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101101; B = 7'b1011110; | Outputs: P=%b | Expected: P=%d",
                 269,
                 
                 P
                 , 
                 
                 10246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100100; B = 7'b1101101; // Expected: {'P': 3924}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100100; B = 7'b1101101; | Outputs: P=%b | Expected: P=%d",
                 270,
                 
                 P
                 , 
                 
                 3924
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101111; B = 7'b1001111; // Expected: {'P': 3713}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101111; B = 7'b1001111; | Outputs: P=%b | Expected: P=%d",
                 271,
                 
                 P
                 , 
                 
                 3713
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110000; B = 7'b1101011; // Expected: {'P': 5136}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110000; B = 7'b1101011; | Outputs: P=%b | Expected: P=%d",
                 272,
                 
                 P
                 , 
                 
                 5136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101100; B = 7'b1111000; // Expected: {'P': 5280}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101100; B = 7'b1111000; | Outputs: P=%b | Expected: P=%d",
                 273,
                 
                 P
                 , 
                 
                 5280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010100; B = 7'b1111111; // Expected: {'P': 2540}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010100; B = 7'b1111111; | Outputs: P=%b | Expected: P=%d",
                 274,
                 
                 P
                 , 
                 
                 2540
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100001; B = 7'b0010111; // Expected: {'P': 759}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100001; B = 7'b0010111; | Outputs: P=%b | Expected: P=%d",
                 275,
                 
                 P
                 , 
                 
                 759
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100100; B = 7'b1110101; // Expected: {'P': 4212}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100100; B = 7'b1110101; | Outputs: P=%b | Expected: P=%d",
                 276,
                 
                 P
                 , 
                 
                 4212
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000111; B = 7'b0011101; // Expected: {'P': 2059}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000111; B = 7'b0011101; | Outputs: P=%b | Expected: P=%d",
                 277,
                 
                 P
                 , 
                 
                 2059
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010110; B = 7'b0000101; // Expected: {'P': 430}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010110; B = 7'b0000101; | Outputs: P=%b | Expected: P=%d",
                 278,
                 
                 P
                 , 
                 
                 430
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001101; B = 7'b0011011; // Expected: {'P': 2079}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001101; B = 7'b0011011; | Outputs: P=%b | Expected: P=%d",
                 279,
                 
                 P
                 , 
                 
                 2079
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110101; B = 7'b0000110; // Expected: {'P': 318}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110101; B = 7'b0000110; | Outputs: P=%b | Expected: P=%d",
                 280,
                 
                 P
                 , 
                 
                 318
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101011; B = 7'b1111111; // Expected: {'P': 5461}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101011; B = 7'b1111111; | Outputs: P=%b | Expected: P=%d",
                 281,
                 
                 P
                 , 
                 
                 5461
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001001; B = 7'b1101110; // Expected: {'P': 8030}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001001; B = 7'b1101110; | Outputs: P=%b | Expected: P=%d",
                 282,
                 
                 P
                 , 
                 
                 8030
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001001; B = 7'b0100111; // Expected: {'P': 2847}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001001; B = 7'b0100111; | Outputs: P=%b | Expected: P=%d",
                 283,
                 
                 P
                 , 
                 
                 2847
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001111; B = 7'b1000111; // Expected: {'P': 1065}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001111; B = 7'b1000111; | Outputs: P=%b | Expected: P=%d",
                 284,
                 
                 P
                 , 
                 
                 1065
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011011; B = 7'b0001000; // Expected: {'P': 728}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011011; B = 7'b0001000; | Outputs: P=%b | Expected: P=%d",
                 285,
                 
                 P
                 , 
                 
                 728
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010001; B = 7'b0110101; // Expected: {'P': 4293}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010001; B = 7'b0110101; | Outputs: P=%b | Expected: P=%d",
                 286,
                 
                 P
                 , 
                 
                 4293
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110111; B = 7'b1101111; // Expected: {'P': 13209}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110111; B = 7'b1101111; | Outputs: P=%b | Expected: P=%d",
                 287,
                 
                 P
                 , 
                 
                 13209
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001000; B = 7'b1001011; // Expected: {'P': 5400}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001000; B = 7'b1001011; | Outputs: P=%b | Expected: P=%d",
                 288,
                 
                 P
                 , 
                 
                 5400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110000; B = 7'b0110001; // Expected: {'P': 2352}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110000; B = 7'b0110001; | Outputs: P=%b | Expected: P=%d",
                 289,
                 
                 P
                 , 
                 
                 2352
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111011; B = 7'b1100000; // Expected: {'P': 11808}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111011; B = 7'b1100000; | Outputs: P=%b | Expected: P=%d",
                 290,
                 
                 P
                 , 
                 
                 11808
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001000; B = 7'b1100010; // Expected: {'P': 784}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001000; B = 7'b1100010; | Outputs: P=%b | Expected: P=%d",
                 291,
                 
                 P
                 , 
                 
                 784
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111111; B = 7'b1110001; // Expected: {'P': 7119}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111111; B = 7'b1110001; | Outputs: P=%b | Expected: P=%d",
                 292,
                 
                 P
                 , 
                 
                 7119
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000111; B = 7'b0011111; // Expected: {'P': 217}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000111; B = 7'b0011111; | Outputs: P=%b | Expected: P=%d",
                 293,
                 
                 P
                 , 
                 
                 217
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011010; B = 7'b1011011; // Expected: {'P': 2366}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011010; B = 7'b1011011; | Outputs: P=%b | Expected: P=%d",
                 294,
                 
                 P
                 , 
                 
                 2366
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110001; B = 7'b0011000; // Expected: {'P': 1176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110001; B = 7'b0011000; | Outputs: P=%b | Expected: P=%d",
                 295,
                 
                 P
                 , 
                 
                 1176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101101; B = 7'b1110100; // Expected: {'P': 5220}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101101; B = 7'b1110100; | Outputs: P=%b | Expected: P=%d",
                 296,
                 
                 P
                 , 
                 
                 5220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001000; B = 7'b0100111; // Expected: {'P': 2808}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001000; B = 7'b0100111; | Outputs: P=%b | Expected: P=%d",
                 297,
                 
                 P
                 , 
                 
                 2808
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010101; B = 7'b0101010; // Expected: {'P': 882}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010101; B = 7'b0101010; | Outputs: P=%b | Expected: P=%d",
                 298,
                 
                 P
                 , 
                 
                 882
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011001; B = 7'b0100100; // Expected: {'P': 3204}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011001; B = 7'b0100100; | Outputs: P=%b | Expected: P=%d",
                 299,
                 
                 P
                 , 
                 
                 3204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110000; B = 7'b0101000; // Expected: {'P': 4480}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110000; B = 7'b0101000; | Outputs: P=%b | Expected: P=%d",
                 300,
                 
                 P
                 , 
                 
                 4480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101001; B = 7'b0101011; // Expected: {'P': 4515}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101001; B = 7'b0101011; | Outputs: P=%b | Expected: P=%d",
                 301,
                 
                 P
                 , 
                 
                 4515
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000000; B = 7'b0010000; // Expected: {'P': 1024}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000000; B = 7'b0010000; | Outputs: P=%b | Expected: P=%d",
                 302,
                 
                 P
                 , 
                 
                 1024
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011001; B = 7'b1100001; // Expected: {'P': 2425}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011001; B = 7'b1100001; | Outputs: P=%b | Expected: P=%d",
                 303,
                 
                 P
                 , 
                 
                 2425
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000011; B = 7'b0111010; // Expected: {'P': 3886}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000011; B = 7'b0111010; | Outputs: P=%b | Expected: P=%d",
                 304,
                 
                 P
                 , 
                 
                 3886
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011001; B = 7'b0101011; // Expected: {'P': 3827}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011001; B = 7'b0101011; | Outputs: P=%b | Expected: P=%d",
                 305,
                 
                 P
                 , 
                 
                 3827
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000101; B = 7'b0000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000101; B = 7'b0000000; | Outputs: P=%b | Expected: P=%d",
                 306,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100101; B = 7'b0110001; // Expected: {'P': 1813}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100101; B = 7'b0110001; | Outputs: P=%b | Expected: P=%d",
                 307,
                 
                 P
                 , 
                 
                 1813
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111001; B = 7'b1010011; // Expected: {'P': 4731}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111001; B = 7'b1010011; | Outputs: P=%b | Expected: P=%d",
                 308,
                 
                 P
                 , 
                 
                 4731
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111111; B = 7'b1110110; // Expected: {'P': 14986}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111111; B = 7'b1110110; | Outputs: P=%b | Expected: P=%d",
                 309,
                 
                 P
                 , 
                 
                 14986
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101010; B = 7'b0111011; // Expected: {'P': 2478}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101010; B = 7'b0111011; | Outputs: P=%b | Expected: P=%d",
                 310,
                 
                 P
                 , 
                 
                 2478
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010011; B = 7'b0111101; // Expected: {'P': 1159}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010011; B = 7'b0111101; | Outputs: P=%b | Expected: P=%d",
                 311,
                 
                 P
                 , 
                 
                 1159
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100101; B = 7'b0100111; // Expected: {'P': 1443}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100101; B = 7'b0100111; | Outputs: P=%b | Expected: P=%d",
                 312,
                 
                 P
                 , 
                 
                 1443
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111011; B = 7'b0000010; // Expected: {'P': 118}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111011; B = 7'b0000010; | Outputs: P=%b | Expected: P=%d",
                 313,
                 
                 P
                 , 
                 
                 118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000110; B = 7'b1000100; // Expected: {'P': 408}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000110; B = 7'b1000100; | Outputs: P=%b | Expected: P=%d",
                 314,
                 
                 P
                 , 
                 
                 408
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101011; B = 7'b1010100; // Expected: {'P': 8988}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101011; B = 7'b1010100; | Outputs: P=%b | Expected: P=%d",
                 315,
                 
                 P
                 , 
                 
                 8988
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101100; B = 7'b0001001; // Expected: {'P': 972}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101100; B = 7'b0001001; | Outputs: P=%b | Expected: P=%d",
                 316,
                 
                 P
                 , 
                 
                 972
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010100; B = 7'b1010001; // Expected: {'P': 1620}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010100; B = 7'b1010001; | Outputs: P=%b | Expected: P=%d",
                 317,
                 
                 P
                 , 
                 
                 1620
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001001; B = 7'b0110110; // Expected: {'P': 486}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001001; B = 7'b0110110; | Outputs: P=%b | Expected: P=%d",
                 318,
                 
                 P
                 , 
                 
                 486
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111101; B = 7'b0000100; // Expected: {'P': 500}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111101; B = 7'b0000100; | Outputs: P=%b | Expected: P=%d",
                 319,
                 
                 P
                 , 
                 
                 500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010010; B = 7'b0011010; // Expected: {'P': 2132}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010010; B = 7'b0011010; | Outputs: P=%b | Expected: P=%d",
                 320,
                 
                 P
                 , 
                 
                 2132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000110; B = 7'b1011111; // Expected: {'P': 570}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000110; B = 7'b1011111; | Outputs: P=%b | Expected: P=%d",
                 321,
                 
                 P
                 , 
                 
                 570
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010111; B = 7'b1000101; // Expected: {'P': 6003}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010111; B = 7'b1000101; | Outputs: P=%b | Expected: P=%d",
                 322,
                 
                 P
                 , 
                 
                 6003
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000001; B = 7'b1011000; // Expected: {'P': 88}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000001; B = 7'b1011000; | Outputs: P=%b | Expected: P=%d",
                 323,
                 
                 P
                 , 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111001; B = 7'b0010010; // Expected: {'P': 2178}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111001; B = 7'b0010010; | Outputs: P=%b | Expected: P=%d",
                 324,
                 
                 P
                 , 
                 
                 2178
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011000; B = 7'b1011001; // Expected: {'P': 7832}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011000; B = 7'b1011001; | Outputs: P=%b | Expected: P=%d",
                 325,
                 
                 P
                 , 
                 
                 7832
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111001; B = 7'b0011111; // Expected: {'P': 1767}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111001; B = 7'b0011111; | Outputs: P=%b | Expected: P=%d",
                 326,
                 
                 P
                 , 
                 
                 1767
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000000; B = 7'b0100101; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000000; B = 7'b0100101; | Outputs: P=%b | Expected: P=%d",
                 327,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110101; B = 7'b0100110; // Expected: {'P': 4446}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110101; B = 7'b0100110; | Outputs: P=%b | Expected: P=%d",
                 328,
                 
                 P
                 , 
                 
                 4446
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101100; B = 7'b1101111; // Expected: {'P': 11988}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101100; B = 7'b1101111; | Outputs: P=%b | Expected: P=%d",
                 329,
                 
                 P
                 , 
                 
                 11988
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011101; B = 7'b1010010; // Expected: {'P': 2378}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011101; B = 7'b1010010; | Outputs: P=%b | Expected: P=%d",
                 330,
                 
                 P
                 , 
                 
                 2378
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111001; B = 7'b1101110; // Expected: {'P': 6270}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111001; B = 7'b1101110; | Outputs: P=%b | Expected: P=%d",
                 331,
                 
                 P
                 , 
                 
                 6270
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000011; B = 7'b1010001; // Expected: {'P': 243}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000011; B = 7'b1010001; | Outputs: P=%b | Expected: P=%d",
                 332,
                 
                 P
                 , 
                 
                 243
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111100; B = 7'b1100001; // Expected: {'P': 12028}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111100; B = 7'b1100001; | Outputs: P=%b | Expected: P=%d",
                 333,
                 
                 P
                 , 
                 
                 12028
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110110; B = 7'b0111100; // Expected: {'P': 7080}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110110; B = 7'b0111100; | Outputs: P=%b | Expected: P=%d",
                 334,
                 
                 P
                 , 
                 
                 7080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011000; B = 7'b1011010; // Expected: {'P': 7920}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011000; B = 7'b1011010; | Outputs: P=%b | Expected: P=%d",
                 335,
                 
                 P
                 , 
                 
                 7920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000010; B = 7'b1100000; // Expected: {'P': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000010; B = 7'b1100000; | Outputs: P=%b | Expected: P=%d",
                 336,
                 
                 P
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000100; B = 7'b1010111; // Expected: {'P': 5916}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000100; B = 7'b1010111; | Outputs: P=%b | Expected: P=%d",
                 337,
                 
                 P
                 , 
                 
                 5916
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011111; B = 7'b1110101; // Expected: {'P': 11115}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011111; B = 7'b1110101; | Outputs: P=%b | Expected: P=%d",
                 338,
                 
                 P
                 , 
                 
                 11115
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101010; B = 7'b0000001; // Expected: {'P': 106}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101010; B = 7'b0000001; | Outputs: P=%b | Expected: P=%d",
                 339,
                 
                 P
                 , 
                 
                 106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100110; B = 7'b1010110; // Expected: {'P': 3268}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100110; B = 7'b1010110; | Outputs: P=%b | Expected: P=%d",
                 340,
                 
                 P
                 , 
                 
                 3268
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111111; B = 7'b0111111; // Expected: {'P': 8001}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111111; B = 7'b0111111; | Outputs: P=%b | Expected: P=%d",
                 341,
                 
                 P
                 , 
                 
                 8001
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010100; B = 7'b0100011; // Expected: {'P': 700}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010100; B = 7'b0100011; | Outputs: P=%b | Expected: P=%d",
                 342,
                 
                 P
                 , 
                 
                 700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100010; B = 7'b0000001; // Expected: {'P': 98}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100010; B = 7'b0000001; | Outputs: P=%b | Expected: P=%d",
                 343,
                 
                 P
                 , 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100100; B = 7'b0000111; // Expected: {'P': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100100; B = 7'b0000111; | Outputs: P=%b | Expected: P=%d",
                 344,
                 
                 P
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001001; B = 7'b1010011; // Expected: {'P': 747}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001001; B = 7'b1010011; | Outputs: P=%b | Expected: P=%d",
                 345,
                 
                 P
                 , 
                 
                 747
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111011; B = 7'b1111111; // Expected: {'P': 7493}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111011; B = 7'b1111111; | Outputs: P=%b | Expected: P=%d",
                 346,
                 
                 P
                 , 
                 
                 7493
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111100; B = 7'b0101100; // Expected: {'P': 5456}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111100; B = 7'b0101100; | Outputs: P=%b | Expected: P=%d",
                 347,
                 
                 P
                 , 
                 
                 5456
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000000; B = 7'b0100010; // Expected: {'P': 2176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000000; B = 7'b0100010; | Outputs: P=%b | Expected: P=%d",
                 348,
                 
                 P
                 , 
                 
                 2176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000001; B = 7'b1000001; // Expected: {'P': 65}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000001; B = 7'b1000001; | Outputs: P=%b | Expected: P=%d",
                 349,
                 
                 P
                 , 
                 
                 65
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110110; B = 7'b0011010; // Expected: {'P': 3068}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110110; B = 7'b0011010; | Outputs: P=%b | Expected: P=%d",
                 350,
                 
                 P
                 , 
                 
                 3068
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010000; B = 7'b0001000; // Expected: {'P': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010000; B = 7'b0001000; | Outputs: P=%b | Expected: P=%d",
                 351,
                 
                 P
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100001; B = 7'b1110001; // Expected: {'P': 10961}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100001; B = 7'b1110001; | Outputs: P=%b | Expected: P=%d",
                 352,
                 
                 P
                 , 
                 
                 10961
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101100; B = 7'b1011101; // Expected: {'P': 10044}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101100; B = 7'b1011101; | Outputs: P=%b | Expected: P=%d",
                 353,
                 
                 P
                 , 
                 
                 10044
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010001; B = 7'b0000001; // Expected: {'P': 81}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010001; B = 7'b0000001; | Outputs: P=%b | Expected: P=%d",
                 354,
                 
                 P
                 , 
                 
                 81
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100010; B = 7'b1110001; // Expected: {'P': 11074}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100010; B = 7'b1110001; | Outputs: P=%b | Expected: P=%d",
                 355,
                 
                 P
                 , 
                 
                 11074
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001111; B = 7'b0111110; // Expected: {'P': 930}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001111; B = 7'b0111110; | Outputs: P=%b | Expected: P=%d",
                 356,
                 
                 P
                 , 
                 
                 930
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111001; B = 7'b0111100; // Expected: {'P': 3420}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111001; B = 7'b0111100; | Outputs: P=%b | Expected: P=%d",
                 357,
                 
                 P
                 , 
                 
                 3420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110001; B = 7'b0101011; // Expected: {'P': 4859}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110001; B = 7'b0101011; | Outputs: P=%b | Expected: P=%d",
                 358,
                 
                 P
                 , 
                 
                 4859
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001101; B = 7'b1000010; // Expected: {'P': 858}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001101; B = 7'b1000010; | Outputs: P=%b | Expected: P=%d",
                 359,
                 
                 P
                 , 
                 
                 858
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011100; B = 7'b1110100; // Expected: {'P': 3248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011100; B = 7'b1110100; | Outputs: P=%b | Expected: P=%d",
                 360,
                 
                 P
                 , 
                 
                 3248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110000; B = 7'b1001000; // Expected: {'P': 3456}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110000; B = 7'b1001000; | Outputs: P=%b | Expected: P=%d",
                 361,
                 
                 P
                 , 
                 
                 3456
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001000; B = 7'b0110100; // Expected: {'P': 416}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001000; B = 7'b0110100; | Outputs: P=%b | Expected: P=%d",
                 362,
                 
                 P
                 , 
                 
                 416
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011110; B = 7'b1010100; // Expected: {'P': 7896}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011110; B = 7'b1010100; | Outputs: P=%b | Expected: P=%d",
                 363,
                 
                 P
                 , 
                 
                 7896
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000000; B = 7'b0011101; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000000; B = 7'b0011101; | Outputs: P=%b | Expected: P=%d",
                 364,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001000; B = 7'b1001101; // Expected: {'P': 616}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001000; B = 7'b1001101; | Outputs: P=%b | Expected: P=%d",
                 365,
                 
                 P
                 , 
                 
                 616
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111010; B = 7'b1010111; // Expected: {'P': 10614}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111010; B = 7'b1010111; | Outputs: P=%b | Expected: P=%d",
                 366,
                 
                 P
                 , 
                 
                 10614
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110011; B = 7'b0000011; // Expected: {'P': 345}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110011; B = 7'b0000011; | Outputs: P=%b | Expected: P=%d",
                 367,
                 
                 P
                 , 
                 
                 345
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010010; B = 7'b0000010; // Expected: {'P': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010010; B = 7'b0000010; | Outputs: P=%b | Expected: P=%d",
                 368,
                 
                 P
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110100; B = 7'b0010111; // Expected: {'P': 1196}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110100; B = 7'b0010111; | Outputs: P=%b | Expected: P=%d",
                 369,
                 
                 P
                 , 
                 
                 1196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111001; B = 7'b0010100; // Expected: {'P': 2420}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111001; B = 7'b0010100; | Outputs: P=%b | Expected: P=%d",
                 370,
                 
                 P
                 , 
                 
                 2420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001101; B = 7'b0101010; // Expected: {'P': 3234}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001101; B = 7'b0101010; | Outputs: P=%b | Expected: P=%d",
                 371,
                 
                 P
                 , 
                 
                 3234
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000010; B = 7'b0010010; // Expected: {'P': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000010; B = 7'b0010010; | Outputs: P=%b | Expected: P=%d",
                 372,
                 
                 P
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000000; B = 7'b0111010; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000000; B = 7'b0111010; | Outputs: P=%b | Expected: P=%d",
                 373,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010101; B = 7'b1111100; // Expected: {'P': 2604}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010101; B = 7'b1111100; | Outputs: P=%b | Expected: P=%d",
                 374,
                 
                 P
                 , 
                 
                 2604
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010010; B = 7'b1100111; // Expected: {'P': 8446}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010010; B = 7'b1100111; | Outputs: P=%b | Expected: P=%d",
                 375,
                 
                 P
                 , 
                 
                 8446
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000010; B = 7'b0111111; // Expected: {'P': 4158}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000010; B = 7'b0111111; | Outputs: P=%b | Expected: P=%d",
                 376,
                 
                 P
                 , 
                 
                 4158
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101110; B = 7'b1111101; // Expected: {'P': 13750}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101110; B = 7'b1111101; | Outputs: P=%b | Expected: P=%d",
                 377,
                 
                 P
                 , 
                 
                 13750
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011011; B = 7'b0100100; // Expected: {'P': 3276}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011011; B = 7'b0100100; | Outputs: P=%b | Expected: P=%d",
                 378,
                 
                 P
                 , 
                 
                 3276
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001110; B = 7'b0001000; // Expected: {'P': 624}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001110; B = 7'b0001000; | Outputs: P=%b | Expected: P=%d",
                 379,
                 
                 P
                 , 
                 
                 624
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110000; B = 7'b1101111; // Expected: {'P': 5328}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110000; B = 7'b1101111; | Outputs: P=%b | Expected: P=%d",
                 380,
                 
                 P
                 , 
                 
                 5328
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110110; B = 7'b1100001; // Expected: {'P': 11446}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110110; B = 7'b1100001; | Outputs: P=%b | Expected: P=%d",
                 381,
                 
                 P
                 , 
                 
                 11446
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111110; B = 7'b1101001; // Expected: {'P': 6510}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111110; B = 7'b1101001; | Outputs: P=%b | Expected: P=%d",
                 382,
                 
                 P
                 , 
                 
                 6510
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010101; B = 7'b1010010; // Expected: {'P': 1722}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010101; B = 7'b1010010; | Outputs: P=%b | Expected: P=%d",
                 383,
                 
                 P
                 , 
                 
                 1722
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011100; B = 7'b1011010; // Expected: {'P': 8280}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011100; B = 7'b1011010; | Outputs: P=%b | Expected: P=%d",
                 384,
                 
                 P
                 , 
                 
                 8280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100011; B = 7'b0110001; // Expected: {'P': 4851}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100011; B = 7'b0110001; | Outputs: P=%b | Expected: P=%d",
                 385,
                 
                 P
                 , 
                 
                 4851
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011110; B = 7'b0111000; // Expected: {'P': 1680}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011110; B = 7'b0111000; | Outputs: P=%b | Expected: P=%d",
                 386,
                 
                 P
                 , 
                 
                 1680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111001; B = 7'b1100011; // Expected: {'P': 11979}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111001; B = 7'b1100011; | Outputs: P=%b | Expected: P=%d",
                 387,
                 
                 P
                 , 
                 
                 11979
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101000; B = 7'b1101000; // Expected: {'P': 10816}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101000; B = 7'b1101000; | Outputs: P=%b | Expected: P=%d",
                 388,
                 
                 P
                 , 
                 
                 10816
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001111; B = 7'b1010011; // Expected: {'P': 1245}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001111; B = 7'b1010011; | Outputs: P=%b | Expected: P=%d",
                 389,
                 
                 P
                 , 
                 
                 1245
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101011; B = 7'b0001000; // Expected: {'P': 856}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101011; B = 7'b0001000; | Outputs: P=%b | Expected: P=%d",
                 390,
                 
                 P
                 , 
                 
                 856
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010010; B = 7'b1101011; // Expected: {'P': 1926}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010010; B = 7'b1101011; | Outputs: P=%b | Expected: P=%d",
                 391,
                 
                 P
                 , 
                 
                 1926
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011011; B = 7'b0111001; // Expected: {'P': 5187}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011011; B = 7'b0111001; | Outputs: P=%b | Expected: P=%d",
                 392,
                 
                 P
                 , 
                 
                 5187
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010101; B = 7'b1100111; // Expected: {'P': 2163}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010101; B = 7'b1100111; | Outputs: P=%b | Expected: P=%d",
                 393,
                 
                 P
                 , 
                 
                 2163
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110111; B = 7'b0011101; // Expected: {'P': 3451}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110111; B = 7'b0011101; | Outputs: P=%b | Expected: P=%d",
                 394,
                 
                 P
                 , 
                 
                 3451
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001011; B = 7'b1110101; // Expected: {'P': 8775}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001011; B = 7'b1110101; | Outputs: P=%b | Expected: P=%d",
                 395,
                 
                 P
                 , 
                 
                 8775
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011110; B = 7'b1001001; // Expected: {'P': 6862}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011110; B = 7'b1001001; | Outputs: P=%b | Expected: P=%d",
                 396,
                 
                 P
                 , 
                 
                 6862
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000110; B = 7'b1101001; // Expected: {'P': 630}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000110; B = 7'b1101001; | Outputs: P=%b | Expected: P=%d",
                 397,
                 
                 P
                 , 
                 
                 630
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110100; B = 7'b0110001; // Expected: {'P': 2548}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110100; B = 7'b0110001; | Outputs: P=%b | Expected: P=%d",
                 398,
                 
                 P
                 , 
                 
                 2548
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000000; B = 7'b1000001; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000000; B = 7'b1000001; | Outputs: P=%b | Expected: P=%d",
                 399,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011111; B = 7'b1111000; // Expected: {'P': 11400}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011111; B = 7'b1111000; | Outputs: P=%b | Expected: P=%d",
                 400,
                 
                 P
                 , 
                 
                 11400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101111; B = 7'b1010100; // Expected: {'P': 3948}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101111; B = 7'b1010100; | Outputs: P=%b | Expected: P=%d",
                 401,
                 
                 P
                 , 
                 
                 3948
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001010; B = 7'b1000000; // Expected: {'P': 4736}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001010; B = 7'b1000000; | Outputs: P=%b | Expected: P=%d",
                 402,
                 
                 P
                 , 
                 
                 4736
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010010; B = 7'b1111010; // Expected: {'P': 2196}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010010; B = 7'b1111010; | Outputs: P=%b | Expected: P=%d",
                 403,
                 
                 P
                 , 
                 
                 2196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101011; B = 7'b0100110; // Expected: {'P': 4066}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101011; B = 7'b0100110; | Outputs: P=%b | Expected: P=%d",
                 404,
                 
                 P
                 , 
                 
                 4066
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001110; B = 7'b0000110; // Expected: {'P': 84}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001110; B = 7'b0000110; | Outputs: P=%b | Expected: P=%d",
                 405,
                 
                 P
                 , 
                 
                 84
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100110; B = 7'b1100111; // Expected: {'P': 10506}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100110; B = 7'b1100111; | Outputs: P=%b | Expected: P=%d",
                 406,
                 
                 P
                 , 
                 
                 10506
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101000; B = 7'b1000000; // Expected: {'P': 2560}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101000; B = 7'b1000000; | Outputs: P=%b | Expected: P=%d",
                 407,
                 
                 P
                 , 
                 
                 2560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001010; B = 7'b0000101; // Expected: {'P': 370}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001010; B = 7'b0000101; | Outputs: P=%b | Expected: P=%d",
                 408,
                 
                 P
                 , 
                 
                 370
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001111; B = 7'b0011001; // Expected: {'P': 1975}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001111; B = 7'b0011001; | Outputs: P=%b | Expected: P=%d",
                 409,
                 
                 P
                 , 
                 
                 1975
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000100; B = 7'b1111001; // Expected: {'P': 8228}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000100; B = 7'b1111001; | Outputs: P=%b | Expected: P=%d",
                 410,
                 
                 P
                 , 
                 
                 8228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100011; B = 7'b1100101; // Expected: {'P': 9999}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100011; B = 7'b1100101; | Outputs: P=%b | Expected: P=%d",
                 411,
                 
                 P
                 , 
                 
                 9999
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001101; B = 7'b1010000; // Expected: {'P': 6160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001101; B = 7'b1010000; | Outputs: P=%b | Expected: P=%d",
                 412,
                 
                 P
                 , 
                 
                 6160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111111; B = 7'b1001000; // Expected: {'P': 9144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111111; B = 7'b1001000; | Outputs: P=%b | Expected: P=%d",
                 413,
                 
                 P
                 , 
                 
                 9144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011010; B = 7'b1101111; // Expected: {'P': 9990}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011010; B = 7'b1101111; | Outputs: P=%b | Expected: P=%d",
                 414,
                 
                 P
                 , 
                 
                 9990
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011010; B = 7'b0101011; // Expected: {'P': 3870}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011010; B = 7'b0101011; | Outputs: P=%b | Expected: P=%d",
                 415,
                 
                 P
                 , 
                 
                 3870
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101001; B = 7'b0010101; // Expected: {'P': 861}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101001; B = 7'b0010101; | Outputs: P=%b | Expected: P=%d",
                 416,
                 
                 P
                 , 
                 
                 861
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111100; B = 7'b1011100; // Expected: {'P': 5520}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111100; B = 7'b1011100; | Outputs: P=%b | Expected: P=%d",
                 417,
                 
                 P
                 , 
                 
                 5520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101001; B = 7'b1011010; // Expected: {'P': 3690}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101001; B = 7'b1011010; | Outputs: P=%b | Expected: P=%d",
                 418,
                 
                 P
                 , 
                 
                 3690
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110011; B = 7'b1100000; // Expected: {'P': 11040}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110011; B = 7'b1100000; | Outputs: P=%b | Expected: P=%d",
                 419,
                 
                 P
                 , 
                 
                 11040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100011; B = 7'b0001101; // Expected: {'P': 455}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100011; B = 7'b0001101; | Outputs: P=%b | Expected: P=%d",
                 420,
                 
                 P
                 , 
                 
                 455
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100110; B = 7'b1000011; // Expected: {'P': 2546}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100110; B = 7'b1000011; | Outputs: P=%b | Expected: P=%d",
                 421,
                 
                 P
                 , 
                 
                 2546
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011110; B = 7'b0101011; // Expected: {'P': 4042}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011110; B = 7'b0101011; | Outputs: P=%b | Expected: P=%d",
                 422,
                 
                 P
                 , 
                 
                 4042
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001101; B = 7'b0011110; // Expected: {'P': 390}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001101; B = 7'b0011110; | Outputs: P=%b | Expected: P=%d",
                 423,
                 
                 P
                 , 
                 
                 390
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000101; B = 7'b1001100; // Expected: {'P': 5244}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000101; B = 7'b1001100; | Outputs: P=%b | Expected: P=%d",
                 424,
                 
                 P
                 , 
                 
                 5244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001110; B = 7'b1111001; // Expected: {'P': 9438}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001110; B = 7'b1111001; | Outputs: P=%b | Expected: P=%d",
                 425,
                 
                 P
                 , 
                 
                 9438
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111101; B = 7'b1011000; // Expected: {'P': 11000}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111101; B = 7'b1011000; | Outputs: P=%b | Expected: P=%d",
                 426,
                 
                 P
                 , 
                 
                 11000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010100; B = 7'b1011110; // Expected: {'P': 1880}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010100; B = 7'b1011110; | Outputs: P=%b | Expected: P=%d",
                 427,
                 
                 P
                 , 
                 
                 1880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000100; B = 7'b1111010; // Expected: {'P': 488}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000100; B = 7'b1111010; | Outputs: P=%b | Expected: P=%d",
                 428,
                 
                 P
                 , 
                 
                 488
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011000; B = 7'b1101110; // Expected: {'P': 9680}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011000; B = 7'b1101110; | Outputs: P=%b | Expected: P=%d",
                 429,
                 
                 P
                 , 
                 
                 9680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010001; B = 7'b1111100; // Expected: {'P': 10044}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010001; B = 7'b1111100; | Outputs: P=%b | Expected: P=%d",
                 430,
                 
                 P
                 , 
                 
                 10044
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101111; B = 7'b0110011; // Expected: {'P': 5661}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101111; B = 7'b0110011; | Outputs: P=%b | Expected: P=%d",
                 431,
                 
                 P
                 , 
                 
                 5661
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010111; B = 7'b0101111; // Expected: {'P': 4089}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010111; B = 7'b0101111; | Outputs: P=%b | Expected: P=%d",
                 432,
                 
                 P
                 , 
                 
                 4089
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100001; B = 7'b1100001; // Expected: {'P': 3201}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100001; B = 7'b1100001; | Outputs: P=%b | Expected: P=%d",
                 433,
                 
                 P
                 , 
                 
                 3201
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010111; B = 7'b0011100; // Expected: {'P': 2436}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010111; B = 7'b0011100; | Outputs: P=%b | Expected: P=%d",
                 434,
                 
                 P
                 , 
                 
                 2436
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011100; B = 7'b0100001; // Expected: {'P': 924}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011100; B = 7'b0100001; | Outputs: P=%b | Expected: P=%d",
                 435,
                 
                 P
                 , 
                 
                 924
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110111; B = 7'b0110010; // Expected: {'P': 2750}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110111; B = 7'b0110010; | Outputs: P=%b | Expected: P=%d",
                 436,
                 
                 P
                 , 
                 
                 2750
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010001; B = 7'b1011001; // Expected: {'P': 1513}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010001; B = 7'b1011001; | Outputs: P=%b | Expected: P=%d",
                 437,
                 
                 P
                 , 
                 
                 1513
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111011; B = 7'b1000101; // Expected: {'P': 4071}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111011; B = 7'b1000101; | Outputs: P=%b | Expected: P=%d",
                 438,
                 
                 P
                 , 
                 
                 4071
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000001; B = 7'b0111001; // Expected: {'P': 57}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000001; B = 7'b0111001; | Outputs: P=%b | Expected: P=%d",
                 439,
                 
                 P
                 , 
                 
                 57
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010011; B = 7'b1001000; // Expected: {'P': 1368}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010011; B = 7'b1001000; | Outputs: P=%b | Expected: P=%d",
                 440,
                 
                 P
                 , 
                 
                 1368
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110001; B = 7'b1110000; // Expected: {'P': 12656}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110001; B = 7'b1110000; | Outputs: P=%b | Expected: P=%d",
                 441,
                 
                 P
                 , 
                 
                 12656
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101101; B = 7'b1011100; // Expected: {'P': 4140}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101101; B = 7'b1011100; | Outputs: P=%b | Expected: P=%d",
                 442,
                 
                 P
                 , 
                 
                 4140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101011; B = 7'b1001110; // Expected: {'P': 3354}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101011; B = 7'b1001110; | Outputs: P=%b | Expected: P=%d",
                 443,
                 
                 P
                 , 
                 
                 3354
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010110; B = 7'b0100011; // Expected: {'P': 3010}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010110; B = 7'b0100011; | Outputs: P=%b | Expected: P=%d",
                 444,
                 
                 P
                 , 
                 
                 3010
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101100; B = 7'b1010110; // Expected: {'P': 3784}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101100; B = 7'b1010110; | Outputs: P=%b | Expected: P=%d",
                 445,
                 
                 P
                 , 
                 
                 3784
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001110; B = 7'b1011010; // Expected: {'P': 1260}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001110; B = 7'b1011010; | Outputs: P=%b | Expected: P=%d",
                 446,
                 
                 P
                 , 
                 
                 1260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110010; B = 7'b1100000; // Expected: {'P': 4800}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110010; B = 7'b1100000; | Outputs: P=%b | Expected: P=%d",
                 447,
                 
                 P
                 , 
                 
                 4800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111011; B = 7'b1111100; // Expected: {'P': 15252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111011; B = 7'b1111100; | Outputs: P=%b | Expected: P=%d",
                 448,
                 
                 P
                 , 
                 
                 15252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010111; B = 7'b0100001; // Expected: {'P': 759}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010111; B = 7'b0100001; | Outputs: P=%b | Expected: P=%d",
                 449,
                 
                 P
                 , 
                 
                 759
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111000; B = 7'b0111011; // Expected: {'P': 7080}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111000; B = 7'b0111011; | Outputs: P=%b | Expected: P=%d",
                 450,
                 
                 P
                 , 
                 
                 7080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001011; B = 7'b0000011; // Expected: {'P': 225}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001011; B = 7'b0000011; | Outputs: P=%b | Expected: P=%d",
                 451,
                 
                 P
                 , 
                 
                 225
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101101; B = 7'b1010111; // Expected: {'P': 9483}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101101; B = 7'b1010111; | Outputs: P=%b | Expected: P=%d",
                 452,
                 
                 P
                 , 
                 
                 9483
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000011; B = 7'b0011000; // Expected: {'P': 1608}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000011; B = 7'b0011000; | Outputs: P=%b | Expected: P=%d",
                 453,
                 
                 P
                 , 
                 
                 1608
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000101; B = 7'b1110001; // Expected: {'P': 565}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000101; B = 7'b1110001; | Outputs: P=%b | Expected: P=%d",
                 454,
                 
                 P
                 , 
                 
                 565
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110110; B = 7'b0111000; // Expected: {'P': 3024}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110110; B = 7'b0111000; | Outputs: P=%b | Expected: P=%d",
                 455,
                 
                 P
                 , 
                 
                 3024
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100000; B = 7'b1001110; // Expected: {'P': 7488}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100000; B = 7'b1001110; | Outputs: P=%b | Expected: P=%d",
                 456,
                 
                 P
                 , 
                 
                 7488
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101100; B = 7'b1101000; // Expected: {'P': 4576}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101100; B = 7'b1101000; | Outputs: P=%b | Expected: P=%d",
                 457,
                 
                 P
                 , 
                 
                 4576
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100000; B = 7'b0001101; // Expected: {'P': 1248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100000; B = 7'b0001101; | Outputs: P=%b | Expected: P=%d",
                 458,
                 
                 P
                 , 
                 
                 1248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101101; B = 7'b1001110; // Expected: {'P': 8502}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101101; B = 7'b1001110; | Outputs: P=%b | Expected: P=%d",
                 459,
                 
                 P
                 , 
                 
                 8502
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110110; B = 7'b0101101; // Expected: {'P': 2430}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110110; B = 7'b0101101; | Outputs: P=%b | Expected: P=%d",
                 460,
                 
                 P
                 , 
                 
                 2430
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011010; B = 7'b1110001; // Expected: {'P': 10170}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011010; B = 7'b1110001; | Outputs: P=%b | Expected: P=%d",
                 461,
                 
                 P
                 , 
                 
                 10170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000100; B = 7'b1100001; // Expected: {'P': 388}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000100; B = 7'b1100001; | Outputs: P=%b | Expected: P=%d",
                 462,
                 
                 P
                 , 
                 
                 388
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000101; B = 7'b0101001; // Expected: {'P': 205}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000101; B = 7'b0101001; | Outputs: P=%b | Expected: P=%d",
                 463,
                 
                 P
                 , 
                 
                 205
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100000; B = 7'b0000001; // Expected: {'P': 32}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100000; B = 7'b0000001; | Outputs: P=%b | Expected: P=%d",
                 464,
                 
                 P
                 , 
                 
                 32
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110010; B = 7'b0100000; // Expected: {'P': 1600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110010; B = 7'b0100000; | Outputs: P=%b | Expected: P=%d",
                 465,
                 
                 P
                 , 
                 
                 1600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101010; B = 7'b1110111; // Expected: {'P': 4998}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101010; B = 7'b1110111; | Outputs: P=%b | Expected: P=%d",
                 466,
                 
                 P
                 , 
                 
                 4998
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010101; B = 7'b0100110; // Expected: {'P': 798}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010101; B = 7'b0100110; | Outputs: P=%b | Expected: P=%d",
                 467,
                 
                 P
                 , 
                 
                 798
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111101; B = 7'b1001100; // Expected: {'P': 4636}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111101; B = 7'b1001100; | Outputs: P=%b | Expected: P=%d",
                 468,
                 
                 P
                 , 
                 
                 4636
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000000; B = 7'b1001100; // Expected: {'P': 4864}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000000; B = 7'b1001100; | Outputs: P=%b | Expected: P=%d",
                 469,
                 
                 P
                 , 
                 
                 4864
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110000; B = 7'b0000101; // Expected: {'P': 560}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110000; B = 7'b0000101; | Outputs: P=%b | Expected: P=%d",
                 470,
                 
                 P
                 , 
                 
                 560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011110; B = 7'b1001111; // Expected: {'P': 2370}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011110; B = 7'b1001111; | Outputs: P=%b | Expected: P=%d",
                 471,
                 
                 P
                 , 
                 
                 2370
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101101; B = 7'b1100000; // Expected: {'P': 10464}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101101; B = 7'b1100000; | Outputs: P=%b | Expected: P=%d",
                 472,
                 
                 P
                 , 
                 
                 10464
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011010; B = 7'b1110000; // Expected: {'P': 2912}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011010; B = 7'b1110000; | Outputs: P=%b | Expected: P=%d",
                 473,
                 
                 P
                 , 
                 
                 2912
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101011; B = 7'b1011101; // Expected: {'P': 3999}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101011; B = 7'b1011101; | Outputs: P=%b | Expected: P=%d",
                 474,
                 
                 P
                 , 
                 
                 3999
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100000; B = 7'b1011110; // Expected: {'P': 3008}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100000; B = 7'b1011110; | Outputs: P=%b | Expected: P=%d",
                 475,
                 
                 P
                 , 
                 
                 3008
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110010; B = 7'b1010000; // Expected: {'P': 9120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110010; B = 7'b1010000; | Outputs: P=%b | Expected: P=%d",
                 476,
                 
                 P
                 , 
                 
                 9120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000001; B = 7'b0011010; // Expected: {'P': 26}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000001; B = 7'b0011010; | Outputs: P=%b | Expected: P=%d",
                 477,
                 
                 P
                 , 
                 
                 26
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101110; B = 7'b0011101; // Expected: {'P': 1334}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101110; B = 7'b0011101; | Outputs: P=%b | Expected: P=%d",
                 478,
                 
                 P
                 , 
                 
                 1334
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000000; B = 7'b1101000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000000; B = 7'b1101000; | Outputs: P=%b | Expected: P=%d",
                 479,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100011; B = 7'b1110111; // Expected: {'P': 4165}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100011; B = 7'b1110111; | Outputs: P=%b | Expected: P=%d",
                 480,
                 
                 P
                 , 
                 
                 4165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111101; B = 7'b0011001; // Expected: {'P': 3125}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111101; B = 7'b0011001; | Outputs: P=%b | Expected: P=%d",
                 481,
                 
                 P
                 , 
                 
                 3125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111001; B = 7'b1011011; // Expected: {'P': 11011}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111001; B = 7'b1011011; | Outputs: P=%b | Expected: P=%d",
                 482,
                 
                 P
                 , 
                 
                 11011
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110000; B = 7'b0110000; // Expected: {'P': 5376}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110000; B = 7'b0110000; | Outputs: P=%b | Expected: P=%d",
                 483,
                 
                 P
                 , 
                 
                 5376
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000110; B = 7'b0110001; // Expected: {'P': 294}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000110; B = 7'b0110001; | Outputs: P=%b | Expected: P=%d",
                 484,
                 
                 P
                 , 
                 
                 294
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011110; B = 7'b1100001; // Expected: {'P': 9118}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011110; B = 7'b1100001; | Outputs: P=%b | Expected: P=%d",
                 485,
                 
                 P
                 , 
                 
                 9118
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010111; B = 7'b0101110; // Expected: {'P': 1058}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010111; B = 7'b0101110; | Outputs: P=%b | Expected: P=%d",
                 486,
                 
                 P
                 , 
                 
                 1058
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110111; B = 7'b0111011; // Expected: {'P': 3245}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110111; B = 7'b0111011; | Outputs: P=%b | Expected: P=%d",
                 487,
                 
                 P
                 , 
                 
                 3245
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110101; B = 7'b1111001; // Expected: {'P': 6413}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110101; B = 7'b1111001; | Outputs: P=%b | Expected: P=%d",
                 488,
                 
                 P
                 , 
                 
                 6413
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010100; B = 7'b0110010; // Expected: {'P': 1000}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010100; B = 7'b0110010; | Outputs: P=%b | Expected: P=%d",
                 489,
                 
                 P
                 , 
                 
                 1000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111001; B = 7'b1101111; // Expected: {'P': 6327}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111001; B = 7'b1101111; | Outputs: P=%b | Expected: P=%d",
                 490,
                 
                 P
                 , 
                 
                 6327
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101100; B = 7'b0111001; // Expected: {'P': 6156}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101100; B = 7'b0111001; | Outputs: P=%b | Expected: P=%d",
                 491,
                 
                 P
                 , 
                 
                 6156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000100; B = 7'b0011101; // Expected: {'P': 116}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000100; B = 7'b0011101; | Outputs: P=%b | Expected: P=%d",
                 492,
                 
                 P
                 , 
                 
                 116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000011; B = 7'b1010010; // Expected: {'P': 246}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000011; B = 7'b1010010; | Outputs: P=%b | Expected: P=%d",
                 493,
                 
                 P
                 , 
                 
                 246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111110; B = 7'b0010100; // Expected: {'P': 2520}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111110; B = 7'b0010100; | Outputs: P=%b | Expected: P=%d",
                 494,
                 
                 P
                 , 
                 
                 2520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001110; B = 7'b1010000; // Expected: {'P': 1120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001110; B = 7'b1010000; | Outputs: P=%b | Expected: P=%d",
                 495,
                 
                 P
                 , 
                 
                 1120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111100; B = 7'b0101111; // Expected: {'P': 5828}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111100; B = 7'b0101111; | Outputs: P=%b | Expected: P=%d",
                 496,
                 
                 P
                 , 
                 
                 5828
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010111; B = 7'b0010011; // Expected: {'P': 1653}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010111; B = 7'b0010011; | Outputs: P=%b | Expected: P=%d",
                 497,
                 
                 P
                 , 
                 
                 1653
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000010; B = 7'b1010111; // Expected: {'P': 5742}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000010; B = 7'b1010111; | Outputs: P=%b | Expected: P=%d",
                 498,
                 
                 P
                 , 
                 
                 5742
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011101; B = 7'b0110100; // Expected: {'P': 4836}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011101; B = 7'b0110100; | Outputs: P=%b | Expected: P=%d",
                 499,
                 
                 P
                 , 
                 
                 4836
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011100; B = 7'b0010010; // Expected: {'P': 1656}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011100; B = 7'b0010010; | Outputs: P=%b | Expected: P=%d",
                 500,
                 
                 P
                 , 
                 
                 1656
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011000; B = 7'b1010001; // Expected: {'P': 1944}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011000; B = 7'b1010001; | Outputs: P=%b | Expected: P=%d",
                 501,
                 
                 P
                 , 
                 
                 1944
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001110; B = 7'b0001110; // Expected: {'P': 1092}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001110; B = 7'b0001110; | Outputs: P=%b | Expected: P=%d",
                 502,
                 
                 P
                 , 
                 
                 1092
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110001; B = 7'b1010001; // Expected: {'P': 3969}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110001; B = 7'b1010001; | Outputs: P=%b | Expected: P=%d",
                 503,
                 
                 P
                 , 
                 
                 3969
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100000; B = 7'b0110000; // Expected: {'P': 4608}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100000; B = 7'b0110000; | Outputs: P=%b | Expected: P=%d",
                 504,
                 
                 P
                 , 
                 
                 4608
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000100; B = 7'b0001000; // Expected: {'P': 544}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000100; B = 7'b0001000; | Outputs: P=%b | Expected: P=%d",
                 505,
                 
                 P
                 , 
                 
                 544
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001000; B = 7'b1001000; // Expected: {'P': 5184}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001000; B = 7'b1001000; | Outputs: P=%b | Expected: P=%d",
                 506,
                 
                 P
                 , 
                 
                 5184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001101; B = 7'b1101110; // Expected: {'P': 8470}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001101; B = 7'b1101110; | Outputs: P=%b | Expected: P=%d",
                 507,
                 
                 P
                 , 
                 
                 8470
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111111; B = 7'b1101111; // Expected: {'P': 6993}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111111; B = 7'b1101111; | Outputs: P=%b | Expected: P=%d",
                 508,
                 
                 P
                 , 
                 
                 6993
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111000; B = 7'b1101010; // Expected: {'P': 5936}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111000; B = 7'b1101010; | Outputs: P=%b | Expected: P=%d",
                 509,
                 
                 P
                 , 
                 
                 5936
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010000; B = 7'b1001110; // Expected: {'P': 1248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010000; B = 7'b1001110; | Outputs: P=%b | Expected: P=%d",
                 510,
                 
                 P
                 , 
                 
                 1248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100011; B = 7'b0011101; // Expected: {'P': 1015}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100011; B = 7'b0011101; | Outputs: P=%b | Expected: P=%d",
                 511,
                 
                 P
                 , 
                 
                 1015
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100011; B = 7'b0011110; // Expected: {'P': 1050}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100011; B = 7'b0011110; | Outputs: P=%b | Expected: P=%d",
                 512,
                 
                 P
                 , 
                 
                 1050
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000011; B = 7'b0001111; // Expected: {'P': 1005}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000011; B = 7'b0001111; | Outputs: P=%b | Expected: P=%d",
                 513,
                 
                 P
                 , 
                 
                 1005
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011011; B = 7'b1101000; // Expected: {'P': 9464}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011011; B = 7'b1101000; | Outputs: P=%b | Expected: P=%d",
                 514,
                 
                 P
                 , 
                 
                 9464
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000100; B = 7'b1110101; // Expected: {'P': 7956}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000100; B = 7'b1110101; | Outputs: P=%b | Expected: P=%d",
                 515,
                 
                 P
                 , 
                 
                 7956
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110011; B = 7'b1110001; // Expected: {'P': 5763}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110011; B = 7'b1110001; | Outputs: P=%b | Expected: P=%d",
                 516,
                 
                 P
                 , 
                 
                 5763
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111101; B = 7'b1000001; // Expected: {'P': 8125}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111101; B = 7'b1000001; | Outputs: P=%b | Expected: P=%d",
                 517,
                 
                 P
                 , 
                 
                 8125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110101; B = 7'b0010110; // Expected: {'P': 2574}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110101; B = 7'b0010110; | Outputs: P=%b | Expected: P=%d",
                 518,
                 
                 P
                 , 
                 
                 2574
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100100; B = 7'b1110100; // Expected: {'P': 4176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100100; B = 7'b1110100; | Outputs: P=%b | Expected: P=%d",
                 519,
                 
                 P
                 , 
                 
                 4176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101001; B = 7'b0110001; // Expected: {'P': 5145}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101001; B = 7'b0110001; | Outputs: P=%b | Expected: P=%d",
                 520,
                 
                 P
                 , 
                 
                 5145
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101000; B = 7'b1000111; // Expected: {'P': 7384}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101000; B = 7'b1000111; | Outputs: P=%b | Expected: P=%d",
                 521,
                 
                 P
                 , 
                 
                 7384
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111110; B = 7'b1101111; // Expected: {'P': 6882}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111110; B = 7'b1101111; | Outputs: P=%b | Expected: P=%d",
                 522,
                 
                 P
                 , 
                 
                 6882
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010111; B = 7'b0000110; // Expected: {'P': 522}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010111; B = 7'b0000110; | Outputs: P=%b | Expected: P=%d",
                 523,
                 
                 P
                 , 
                 
                 522
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001010; B = 7'b1100000; // Expected: {'P': 960}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001010; B = 7'b1100000; | Outputs: P=%b | Expected: P=%d",
                 524,
                 
                 P
                 , 
                 
                 960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101000; B = 7'b0101100; // Expected: {'P': 1760}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101000; B = 7'b0101100; | Outputs: P=%b | Expected: P=%d",
                 525,
                 
                 P
                 , 
                 
                 1760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011111; B = 7'b1101110; // Expected: {'P': 10450}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011111; B = 7'b1101110; | Outputs: P=%b | Expected: P=%d",
                 526,
                 
                 P
                 , 
                 
                 10450
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010101; B = 7'b1101100; // Expected: {'P': 9180}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010101; B = 7'b1101100; | Outputs: P=%b | Expected: P=%d",
                 527,
                 
                 P
                 , 
                 
                 9180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101001; B = 7'b1100001; // Expected: {'P': 10185}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101001; B = 7'b1100001; | Outputs: P=%b | Expected: P=%d",
                 528,
                 
                 P
                 , 
                 
                 10185
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101010; B = 7'b1011111; // Expected: {'P': 3990}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101010; B = 7'b1011111; | Outputs: P=%b | Expected: P=%d",
                 529,
                 
                 P
                 , 
                 
                 3990
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110111; B = 7'b1111011; // Expected: {'P': 6765}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110111; B = 7'b1111011; | Outputs: P=%b | Expected: P=%d",
                 530,
                 
                 P
                 , 
                 
                 6765
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111011; B = 7'b0011110; // Expected: {'P': 3690}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111011; B = 7'b0011110; | Outputs: P=%b | Expected: P=%d",
                 531,
                 
                 P
                 , 
                 
                 3690
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010110; B = 7'b0000110; // Expected: {'P': 132}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010110; B = 7'b0000110; | Outputs: P=%b | Expected: P=%d",
                 532,
                 
                 P
                 , 
                 
                 132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000010; B = 7'b0010010; // Expected: {'P': 1188}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000010; B = 7'b0010010; | Outputs: P=%b | Expected: P=%d",
                 533,
                 
                 P
                 , 
                 
                 1188
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001110; B = 7'b0011001; // Expected: {'P': 1950}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001110; B = 7'b0011001; | Outputs: P=%b | Expected: P=%d",
                 534,
                 
                 P
                 , 
                 
                 1950
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000001; B = 7'b0010010; // Expected: {'P': 1170}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000001; B = 7'b0010010; | Outputs: P=%b | Expected: P=%d",
                 535,
                 
                 P
                 , 
                 
                 1170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101011; B = 7'b0100111; // Expected: {'P': 4173}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101011; B = 7'b0100111; | Outputs: P=%b | Expected: P=%d",
                 536,
                 
                 P
                 , 
                 
                 4173
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011111; B = 7'b1100101; // Expected: {'P': 3131}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011111; B = 7'b1100101; | Outputs: P=%b | Expected: P=%d",
                 537,
                 
                 P
                 , 
                 
                 3131
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110010; B = 7'b0000010; // Expected: {'P': 100}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110010; B = 7'b0000010; | Outputs: P=%b | Expected: P=%d",
                 538,
                 
                 P
                 , 
                 
                 100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111100; B = 7'b0000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111100; B = 7'b0000000; | Outputs: P=%b | Expected: P=%d",
                 539,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011100; B = 7'b0010011; // Expected: {'P': 1748}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011100; B = 7'b0010011; | Outputs: P=%b | Expected: P=%d",
                 540,
                 
                 P
                 , 
                 
                 1748
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000011; B = 7'b0000110; // Expected: {'P': 18}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000011; B = 7'b0000110; | Outputs: P=%b | Expected: P=%d",
                 541,
                 
                 P
                 , 
                 
                 18
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100101; B = 7'b0111010; // Expected: {'P': 2146}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100101; B = 7'b0111010; | Outputs: P=%b | Expected: P=%d",
                 542,
                 
                 P
                 , 
                 
                 2146
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111100; B = 7'b1111010; // Expected: {'P': 15128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111100; B = 7'b1111010; | Outputs: P=%b | Expected: P=%d",
                 543,
                 
                 P
                 , 
                 
                 15128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001000; B = 7'b0110000; // Expected: {'P': 384}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001000; B = 7'b0110000; | Outputs: P=%b | Expected: P=%d",
                 544,
                 
                 P
                 , 
                 
                 384
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101001; B = 7'b1000000; // Expected: {'P': 2624}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101001; B = 7'b1000000; | Outputs: P=%b | Expected: P=%d",
                 545,
                 
                 P
                 , 
                 
                 2624
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000100; B = 7'b1011111; // Expected: {'P': 380}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000100; B = 7'b1011111; | Outputs: P=%b | Expected: P=%d",
                 546,
                 
                 P
                 , 
                 
                 380
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100110; B = 7'b1100111; // Expected: {'P': 3914}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100110; B = 7'b1100111; | Outputs: P=%b | Expected: P=%d",
                 547,
                 
                 P
                 , 
                 
                 3914
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000001; B = 7'b0111100; // Expected: {'P': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000001; B = 7'b0111100; | Outputs: P=%b | Expected: P=%d",
                 548,
                 
                 P
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010001; B = 7'b0110010; // Expected: {'P': 850}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010001; B = 7'b0110010; | Outputs: P=%b | Expected: P=%d",
                 549,
                 
                 P
                 , 
                 
                 850
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111011; B = 7'b0100110; // Expected: {'P': 4674}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111011; B = 7'b0100110; | Outputs: P=%b | Expected: P=%d",
                 550,
                 
                 P
                 , 
                 
                 4674
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001001; B = 7'b0110010; // Expected: {'P': 3650}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001001; B = 7'b0110010; | Outputs: P=%b | Expected: P=%d",
                 551,
                 
                 P
                 , 
                 
                 3650
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100100; B = 7'b0101101; // Expected: {'P': 1620}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100100; B = 7'b0101101; | Outputs: P=%b | Expected: P=%d",
                 552,
                 
                 P
                 , 
                 
                 1620
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110111; B = 7'b0100101; // Expected: {'P': 4403}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110111; B = 7'b0100101; | Outputs: P=%b | Expected: P=%d",
                 553,
                 
                 P
                 , 
                 
                 4403
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000100; B = 7'b0110000; // Expected: {'P': 3264}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000100; B = 7'b0110000; | Outputs: P=%b | Expected: P=%d",
                 554,
                 
                 P
                 , 
                 
                 3264
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011001; B = 7'b1000100; // Expected: {'P': 1700}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011001; B = 7'b1000100; | Outputs: P=%b | Expected: P=%d",
                 555,
                 
                 P
                 , 
                 
                 1700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101110; B = 7'b0001101; // Expected: {'P': 1430}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101110; B = 7'b0001101; | Outputs: P=%b | Expected: P=%d",
                 556,
                 
                 P
                 , 
                 
                 1430
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100101; B = 7'b0100001; // Expected: {'P': 1221}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100101; B = 7'b0100001; | Outputs: P=%b | Expected: P=%d",
                 557,
                 
                 P
                 , 
                 
                 1221
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010000; B = 7'b0001001; // Expected: {'P': 720}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010000; B = 7'b0001001; | Outputs: P=%b | Expected: P=%d",
                 558,
                 
                 P
                 , 
                 
                 720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010110; B = 7'b0101011; // Expected: {'P': 3698}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010110; B = 7'b0101011; | Outputs: P=%b | Expected: P=%d",
                 559,
                 
                 P
                 , 
                 
                 3698
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111110; B = 7'b1000001; // Expected: {'P': 8190}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111110; B = 7'b1000001; | Outputs: P=%b | Expected: P=%d",
                 560,
                 
                 P
                 , 
                 
                 8190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010100; B = 7'b1110111; // Expected: {'P': 9996}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010100; B = 7'b1110111; | Outputs: P=%b | Expected: P=%d",
                 561,
                 
                 P
                 , 
                 
                 9996
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001100; B = 7'b0001110; // Expected: {'P': 1064}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001100; B = 7'b0001110; | Outputs: P=%b | Expected: P=%d",
                 562,
                 
                 P
                 , 
                 
                 1064
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001110; B = 7'b0010000; // Expected: {'P': 1248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001110; B = 7'b0010000; | Outputs: P=%b | Expected: P=%d",
                 563,
                 
                 P
                 , 
                 
                 1248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010100; B = 7'b1001001; // Expected: {'P': 1460}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010100; B = 7'b1001001; | Outputs: P=%b | Expected: P=%d",
                 564,
                 
                 P
                 , 
                 
                 1460
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111001; B = 7'b0110110; // Expected: {'P': 3078}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111001; B = 7'b0110110; | Outputs: P=%b | Expected: P=%d",
                 565,
                 
                 P
                 , 
                 
                 3078
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001011; B = 7'b1100011; // Expected: {'P': 1089}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001011; B = 7'b1100011; | Outputs: P=%b | Expected: P=%d",
                 566,
                 
                 P
                 , 
                 
                 1089
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000000; B = 7'b1111100; // Expected: {'P': 7936}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000000; B = 7'b1111100; | Outputs: P=%b | Expected: P=%d",
                 567,
                 
                 P
                 , 
                 
                 7936
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101100; B = 7'b1100000; // Expected: {'P': 10368}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101100; B = 7'b1100000; | Outputs: P=%b | Expected: P=%d",
                 568,
                 
                 P
                 , 
                 
                 10368
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100100; B = 7'b0101010; // Expected: {'P': 4200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100100; B = 7'b0101010; | Outputs: P=%b | Expected: P=%d",
                 569,
                 
                 P
                 , 
                 
                 4200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010110; B = 7'b1000010; // Expected: {'P': 5676}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010110; B = 7'b1000010; | Outputs: P=%b | Expected: P=%d",
                 570,
                 
                 P
                 , 
                 
                 5676
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100101; B = 7'b0000011; // Expected: {'P': 111}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100101; B = 7'b0000011; | Outputs: P=%b | Expected: P=%d",
                 571,
                 
                 P
                 , 
                 
                 111
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010011; B = 7'b0001100; // Expected: {'P': 228}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010011; B = 7'b0001100; | Outputs: P=%b | Expected: P=%d",
                 572,
                 
                 P
                 , 
                 
                 228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110101; B = 7'b1100000; // Expected: {'P': 11232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110101; B = 7'b1100000; | Outputs: P=%b | Expected: P=%d",
                 573,
                 
                 P
                 , 
                 
                 11232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011011; B = 7'b1011110; // Expected: {'P': 2538}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011011; B = 7'b1011110; | Outputs: P=%b | Expected: P=%d",
                 574,
                 
                 P
                 , 
                 
                 2538
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111110; B = 7'b1001111; // Expected: {'P': 4898}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111110; B = 7'b1001111; | Outputs: P=%b | Expected: P=%d",
                 575,
                 
                 P
                 , 
                 
                 4898
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111001; B = 7'b0000110; // Expected: {'P': 342}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111001; B = 7'b0000110; | Outputs: P=%b | Expected: P=%d",
                 576,
                 
                 P
                 , 
                 
                 342
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000101; B = 7'b1100110; // Expected: {'P': 510}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000101; B = 7'b1100110; | Outputs: P=%b | Expected: P=%d",
                 577,
                 
                 P
                 , 
                 
                 510
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101011; B = 7'b1100101; // Expected: {'P': 4343}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101011; B = 7'b1100101; | Outputs: P=%b | Expected: P=%d",
                 578,
                 
                 P
                 , 
                 
                 4343
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011011; B = 7'b1011010; // Expected: {'P': 8190}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011011; B = 7'b1011010; | Outputs: P=%b | Expected: P=%d",
                 579,
                 
                 P
                 , 
                 
                 8190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100010; B = 7'b1100101; // Expected: {'P': 9898}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100010; B = 7'b1100101; | Outputs: P=%b | Expected: P=%d",
                 580,
                 
                 P
                 , 
                 
                 9898
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100001; B = 7'b1110101; // Expected: {'P': 11349}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100001; B = 7'b1110101; | Outputs: P=%b | Expected: P=%d",
                 581,
                 
                 P
                 , 
                 
                 11349
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011000; B = 7'b0101110; // Expected: {'P': 4048}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011000; B = 7'b0101110; | Outputs: P=%b | Expected: P=%d",
                 582,
                 
                 P
                 , 
                 
                 4048
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101001; B = 7'b0000111; // Expected: {'P': 735}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101001; B = 7'b0000111; | Outputs: P=%b | Expected: P=%d",
                 583,
                 
                 P
                 , 
                 
                 735
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011011; B = 7'b1101011; // Expected: {'P': 9737}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011011; B = 7'b1101011; | Outputs: P=%b | Expected: P=%d",
                 584,
                 
                 P
                 , 
                 
                 9737
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100010; B = 7'b1111101; // Expected: {'P': 12250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100010; B = 7'b1111101; | Outputs: P=%b | Expected: P=%d",
                 585,
                 
                 P
                 , 
                 
                 12250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000011; B = 7'b1100100; // Expected: {'P': 300}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000011; B = 7'b1100100; | Outputs: P=%b | Expected: P=%d",
                 586,
                 
                 P
                 , 
                 
                 300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100000; B = 7'b0111000; // Expected: {'P': 1792}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100000; B = 7'b0111000; | Outputs: P=%b | Expected: P=%d",
                 587,
                 
                 P
                 , 
                 
                 1792
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011111; B = 7'b0111001; // Expected: {'P': 1767}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011111; B = 7'b0111001; | Outputs: P=%b | Expected: P=%d",
                 588,
                 
                 P
                 , 
                 
                 1767
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010100; B = 7'b1011100; // Expected: {'P': 1840}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010100; B = 7'b1011100; | Outputs: P=%b | Expected: P=%d",
                 589,
                 
                 P
                 , 
                 
                 1840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110011; B = 7'b0111001; // Expected: {'P': 2907}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110011; B = 7'b0111001; | Outputs: P=%b | Expected: P=%d",
                 590,
                 
                 P
                 , 
                 
                 2907
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100000; B = 7'b1100111; // Expected: {'P': 9888}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100000; B = 7'b1100111; | Outputs: P=%b | Expected: P=%d",
                 591,
                 
                 P
                 , 
                 
                 9888
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011011; B = 7'b0011100; // Expected: {'P': 2548}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011011; B = 7'b0011100; | Outputs: P=%b | Expected: P=%d",
                 592,
                 
                 P
                 , 
                 
                 2548
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000100; B = 7'b1101100; // Expected: {'P': 7344}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000100; B = 7'b1101100; | Outputs: P=%b | Expected: P=%d",
                 593,
                 
                 P
                 , 
                 
                 7344
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111001; B = 7'b0100010; // Expected: {'P': 4114}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111001; B = 7'b0100010; | Outputs: P=%b | Expected: P=%d",
                 594,
                 
                 P
                 , 
                 
                 4114
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110000; B = 7'b0011110; // Expected: {'P': 1440}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110000; B = 7'b0011110; | Outputs: P=%b | Expected: P=%d",
                 595,
                 
                 P
                 , 
                 
                 1440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011100; B = 7'b1000110; // Expected: {'P': 6440}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011100; B = 7'b1000110; | Outputs: P=%b | Expected: P=%d",
                 596,
                 
                 P
                 , 
                 
                 6440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001000; B = 7'b1100110; // Expected: {'P': 7344}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001000; B = 7'b1100110; | Outputs: P=%b | Expected: P=%d",
                 597,
                 
                 P
                 , 
                 
                 7344
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111000; B = 7'b0110110; // Expected: {'P': 6480}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111000; B = 7'b0110110; | Outputs: P=%b | Expected: P=%d",
                 598,
                 
                 P
                 , 
                 
                 6480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100111; B = 7'b0011000; // Expected: {'P': 936}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100111; B = 7'b0011000; | Outputs: P=%b | Expected: P=%d",
                 599,
                 
                 P
                 , 
                 
                 936
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100101; B = 7'b1001110; // Expected: {'P': 2886}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100101; B = 7'b1001110; | Outputs: P=%b | Expected: P=%d",
                 600,
                 
                 P
                 , 
                 
                 2886
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010101; B = 7'b1011000; // Expected: {'P': 1848}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010101; B = 7'b1011000; | Outputs: P=%b | Expected: P=%d",
                 601,
                 
                 P
                 , 
                 
                 1848
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100110; B = 7'b0001001; // Expected: {'P': 918}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100110; B = 7'b0001001; | Outputs: P=%b | Expected: P=%d",
                 602,
                 
                 P
                 , 
                 
                 918
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000010; B = 7'b0100111; // Expected: {'P': 78}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000010; B = 7'b0100111; | Outputs: P=%b | Expected: P=%d",
                 603,
                 
                 P
                 , 
                 
                 78
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011111; B = 7'b1011001; // Expected: {'P': 8455}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011111; B = 7'b1011001; | Outputs: P=%b | Expected: P=%d",
                 604,
                 
                 P
                 , 
                 
                 8455
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100001; B = 7'b0111101; // Expected: {'P': 5917}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100001; B = 7'b0111101; | Outputs: P=%b | Expected: P=%d",
                 605,
                 
                 P
                 , 
                 
                 5917
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011010; B = 7'b1010000; // Expected: {'P': 2080}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011010; B = 7'b1010000; | Outputs: P=%b | Expected: P=%d",
                 606,
                 
                 P
                 , 
                 
                 2080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111001; B = 7'b0111000; // Expected: {'P': 6776}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111001; B = 7'b0111000; | Outputs: P=%b | Expected: P=%d",
                 607,
                 
                 P
                 , 
                 
                 6776
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111111; B = 7'b0110011; // Expected: {'P': 6477}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111111; B = 7'b0110011; | Outputs: P=%b | Expected: P=%d",
                 608,
                 
                 P
                 , 
                 
                 6477
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010110; B = 7'b1011011; // Expected: {'P': 7826}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010110; B = 7'b1011011; | Outputs: P=%b | Expected: P=%d",
                 609,
                 
                 P
                 , 
                 
                 7826
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001100; B = 7'b1000101; // Expected: {'P': 828}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001100; B = 7'b1000101; | Outputs: P=%b | Expected: P=%d",
                 610,
                 
                 P
                 , 
                 
                 828
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001101; B = 7'b1110110; // Expected: {'P': 9086}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001101; B = 7'b1110110; | Outputs: P=%b | Expected: P=%d",
                 611,
                 
                 P
                 , 
                 
                 9086
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100010; B = 7'b0001001; // Expected: {'P': 306}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100010; B = 7'b0001001; | Outputs: P=%b | Expected: P=%d",
                 612,
                 
                 P
                 , 
                 
                 306
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011111; B = 7'b1000111; // Expected: {'P': 6745}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011111; B = 7'b1000111; | Outputs: P=%b | Expected: P=%d",
                 613,
                 
                 P
                 , 
                 
                 6745
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110001; B = 7'b1110100; // Expected: {'P': 5684}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110001; B = 7'b1110100; | Outputs: P=%b | Expected: P=%d",
                 614,
                 
                 P
                 , 
                 
                 5684
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011101; B = 7'b1101111; // Expected: {'P': 3219}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011101; B = 7'b1101111; | Outputs: P=%b | Expected: P=%d",
                 615,
                 
                 P
                 , 
                 
                 3219
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111010; B = 7'b0111010; // Expected: {'P': 3364}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111010; B = 7'b0111010; | Outputs: P=%b | Expected: P=%d",
                 616,
                 
                 P
                 , 
                 
                 3364
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010101; B = 7'b0010110; // Expected: {'P': 462}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010101; B = 7'b0010110; | Outputs: P=%b | Expected: P=%d",
                 617,
                 
                 P
                 , 
                 
                 462
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010010; B = 7'b0110100; // Expected: {'P': 936}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010010; B = 7'b0110100; | Outputs: P=%b | Expected: P=%d",
                 618,
                 
                 P
                 , 
                 
                 936
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011111; B = 7'b1101010; // Expected: {'P': 10070}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011111; B = 7'b1101010; | Outputs: P=%b | Expected: P=%d",
                 619,
                 
                 P
                 , 
                 
                 10070
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000110; B = 7'b0110100; // Expected: {'P': 3640}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000110; B = 7'b0110100; | Outputs: P=%b | Expected: P=%d",
                 620,
                 
                 P
                 , 
                 
                 3640
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111011; B = 7'b1000001; // Expected: {'P': 3835}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111011; B = 7'b1000001; | Outputs: P=%b | Expected: P=%d",
                 621,
                 
                 P
                 , 
                 
                 3835
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110101; B = 7'b1101100; // Expected: {'P': 5724}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110101; B = 7'b1101100; | Outputs: P=%b | Expected: P=%d",
                 622,
                 
                 P
                 , 
                 
                 5724
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010011; B = 7'b1000100; // Expected: {'P': 5644}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010011; B = 7'b1000100; | Outputs: P=%b | Expected: P=%d",
                 623,
                 
                 P
                 , 
                 
                 5644
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000111; B = 7'b1100001; // Expected: {'P': 679}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000111; B = 7'b1100001; | Outputs: P=%b | Expected: P=%d",
                 624,
                 
                 P
                 , 
                 
                 679
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111001; B = 7'b1011010; // Expected: {'P': 10890}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111001; B = 7'b1011010; | Outputs: P=%b | Expected: P=%d",
                 625,
                 
                 P
                 , 
                 
                 10890
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111110; B = 7'b0100110; // Expected: {'P': 4788}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111110; B = 7'b0100110; | Outputs: P=%b | Expected: P=%d",
                 626,
                 
                 P
                 , 
                 
                 4788
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001100; B = 7'b1000111; // Expected: {'P': 852}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001100; B = 7'b1000111; | Outputs: P=%b | Expected: P=%d",
                 627,
                 
                 P
                 , 
                 
                 852
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110010; B = 7'b1011110; // Expected: {'P': 4700}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110010; B = 7'b1011110; | Outputs: P=%b | Expected: P=%d",
                 628,
                 
                 P
                 , 
                 
                 4700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001010; B = 7'b0001111; // Expected: {'P': 1110}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001010; B = 7'b0001111; | Outputs: P=%b | Expected: P=%d",
                 629,
                 
                 P
                 , 
                 
                 1110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011101; B = 7'b0000001; // Expected: {'P': 93}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011101; B = 7'b0000001; | Outputs: P=%b | Expected: P=%d",
                 630,
                 
                 P
                 , 
                 
                 93
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010010; B = 7'b0101110; // Expected: {'P': 828}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010010; B = 7'b0101110; | Outputs: P=%b | Expected: P=%d",
                 631,
                 
                 P
                 , 
                 
                 828
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101010; B = 7'b0010101; // Expected: {'P': 2226}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101010; B = 7'b0010101; | Outputs: P=%b | Expected: P=%d",
                 632,
                 
                 P
                 , 
                 
                 2226
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101110; B = 7'b1000000; // Expected: {'P': 2944}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101110; B = 7'b1000000; | Outputs: P=%b | Expected: P=%d",
                 633,
                 
                 P
                 , 
                 
                 2944
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001100; B = 7'b0011000; // Expected: {'P': 288}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001100; B = 7'b0011000; | Outputs: P=%b | Expected: P=%d",
                 634,
                 
                 P
                 , 
                 
                 288
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000000; B = 7'b0111111; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000000; B = 7'b0111111; | Outputs: P=%b | Expected: P=%d",
                 635,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111110; B = 7'b0111010; // Expected: {'P': 7308}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111110; B = 7'b0111010; | Outputs: P=%b | Expected: P=%d",
                 636,
                 
                 P
                 , 
                 
                 7308
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010000; B = 7'b0010010; // Expected: {'P': 1440}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010000; B = 7'b0010010; | Outputs: P=%b | Expected: P=%d",
                 637,
                 
                 P
                 , 
                 
                 1440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010010; B = 7'b0010000; // Expected: {'P': 1312}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010010; B = 7'b0010000; | Outputs: P=%b | Expected: P=%d",
                 638,
                 
                 P
                 , 
                 
                 1312
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111110; B = 7'b1010000; // Expected: {'P': 4960}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111110; B = 7'b1010000; | Outputs: P=%b | Expected: P=%d",
                 639,
                 
                 P
                 , 
                 
                 4960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100010; B = 7'b1000000; // Expected: {'P': 2176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100010; B = 7'b1000000; | Outputs: P=%b | Expected: P=%d",
                 640,
                 
                 P
                 , 
                 
                 2176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110100; B = 7'b0010000; // Expected: {'P': 1856}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110100; B = 7'b0010000; | Outputs: P=%b | Expected: P=%d",
                 641,
                 
                 P
                 , 
                 
                 1856
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111100; B = 7'b1101100; // Expected: {'P': 6480}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111100; B = 7'b1101100; | Outputs: P=%b | Expected: P=%d",
                 642,
                 
                 P
                 , 
                 
                 6480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010110; B = 7'b1000011; // Expected: {'P': 5762}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010110; B = 7'b1000011; | Outputs: P=%b | Expected: P=%d",
                 643,
                 
                 P
                 , 
                 
                 5762
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010101; B = 7'b0100010; // Expected: {'P': 2890}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010101; B = 7'b0100010; | Outputs: P=%b | Expected: P=%d",
                 644,
                 
                 P
                 , 
                 
                 2890
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011101; B = 7'b1101100; // Expected: {'P': 3132}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011101; B = 7'b1101100; | Outputs: P=%b | Expected: P=%d",
                 645,
                 
                 P
                 , 
                 
                 3132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110001; B = 7'b0100010; // Expected: {'P': 3842}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110001; B = 7'b0100010; | Outputs: P=%b | Expected: P=%d",
                 646,
                 
                 P
                 , 
                 
                 3842
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101101; B = 7'b1000001; // Expected: {'P': 7085}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101101; B = 7'b1000001; | Outputs: P=%b | Expected: P=%d",
                 647,
                 
                 P
                 , 
                 
                 7085
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011011; B = 7'b1011001; // Expected: {'P': 2403}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011011; B = 7'b1011001; | Outputs: P=%b | Expected: P=%d",
                 648,
                 
                 P
                 , 
                 
                 2403
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100000; B = 7'b1101010; // Expected: {'P': 3392}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100000; B = 7'b1101010; | Outputs: P=%b | Expected: P=%d",
                 649,
                 
                 P
                 , 
                 
                 3392
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001111; B = 7'b0010101; // Expected: {'P': 1659}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001111; B = 7'b0010101; | Outputs: P=%b | Expected: P=%d",
                 650,
                 
                 P
                 , 
                 
                 1659
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000001; B = 7'b0101101; // Expected: {'P': 2925}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000001; B = 7'b0101101; | Outputs: P=%b | Expected: P=%d",
                 651,
                 
                 P
                 , 
                 
                 2925
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100000; B = 7'b0001001; // Expected: {'P': 288}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100000; B = 7'b0001001; | Outputs: P=%b | Expected: P=%d",
                 652,
                 
                 P
                 , 
                 
                 288
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111111; B = 7'b0110001; // Expected: {'P': 3087}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111111; B = 7'b0110001; | Outputs: P=%b | Expected: P=%d",
                 653,
                 
                 P
                 , 
                 
                 3087
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110010; B = 7'b1101001; // Expected: {'P': 11970}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110010; B = 7'b1101001; | Outputs: P=%b | Expected: P=%d",
                 654,
                 
                 P
                 , 
                 
                 11970
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110010; B = 7'b0000010; // Expected: {'P': 228}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110010; B = 7'b0000010; | Outputs: P=%b | Expected: P=%d",
                 655,
                 
                 P
                 , 
                 
                 228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011111; B = 7'b0011110; // Expected: {'P': 2850}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011111; B = 7'b0011110; | Outputs: P=%b | Expected: P=%d",
                 656,
                 
                 P
                 , 
                 
                 2850
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011011; B = 7'b1101011; // Expected: {'P': 2889}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011011; B = 7'b1101011; | Outputs: P=%b | Expected: P=%d",
                 657,
                 
                 P
                 , 
                 
                 2889
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011000; B = 7'b0101011; // Expected: {'P': 1032}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011000; B = 7'b0101011; | Outputs: P=%b | Expected: P=%d",
                 658,
                 
                 P
                 , 
                 
                 1032
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100010; B = 7'b0111010; // Expected: {'P': 1972}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100010; B = 7'b0111010; | Outputs: P=%b | Expected: P=%d",
                 659,
                 
                 P
                 , 
                 
                 1972
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010000; B = 7'b1110110; // Expected: {'P': 1888}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010000; B = 7'b1110110; | Outputs: P=%b | Expected: P=%d",
                 660,
                 
                 P
                 , 
                 
                 1888
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100111; B = 7'b0000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100111; B = 7'b0000000; | Outputs: P=%b | Expected: P=%d",
                 661,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011000; B = 7'b0001000; // Expected: {'P': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011000; B = 7'b0001000; | Outputs: P=%b | Expected: P=%d",
                 662,
                 
                 P
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001011; B = 7'b0100100; // Expected: {'P': 396}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001011; B = 7'b0100100; | Outputs: P=%b | Expected: P=%d",
                 663,
                 
                 P
                 , 
                 
                 396
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111001; B = 7'b0111001; // Expected: {'P': 3249}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111001; B = 7'b0111001; | Outputs: P=%b | Expected: P=%d",
                 664,
                 
                 P
                 , 
                 
                 3249
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010001; B = 7'b0001011; // Expected: {'P': 187}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010001; B = 7'b0001011; | Outputs: P=%b | Expected: P=%d",
                 665,
                 
                 P
                 , 
                 
                 187
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111101; B = 7'b1011000; // Expected: {'P': 5368}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111101; B = 7'b1011000; | Outputs: P=%b | Expected: P=%d",
                 666,
                 
                 P
                 , 
                 
                 5368
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101001; B = 7'b0000101; // Expected: {'P': 525}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101001; B = 7'b0000101; | Outputs: P=%b | Expected: P=%d",
                 667,
                 
                 P
                 , 
                 
                 525
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010000; B = 7'b0101010; // Expected: {'P': 672}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010000; B = 7'b0101010; | Outputs: P=%b | Expected: P=%d",
                 668,
                 
                 P
                 , 
                 
                 672
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001010; B = 7'b0101011; // Expected: {'P': 3182}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001010; B = 7'b0101011; | Outputs: P=%b | Expected: P=%d",
                 669,
                 
                 P
                 , 
                 
                 3182
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110111; B = 7'b0011110; // Expected: {'P': 3570}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110111; B = 7'b0011110; | Outputs: P=%b | Expected: P=%d",
                 670,
                 
                 P
                 , 
                 
                 3570
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100010; B = 7'b0011011; // Expected: {'P': 918}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100010; B = 7'b0011011; | Outputs: P=%b | Expected: P=%d",
                 671,
                 
                 P
                 , 
                 
                 918
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011101; B = 7'b0011000; // Expected: {'P': 2232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011101; B = 7'b0011000; | Outputs: P=%b | Expected: P=%d",
                 672,
                 
                 P
                 , 
                 
                 2232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011111; B = 7'b0011001; // Expected: {'P': 2375}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011111; B = 7'b0011001; | Outputs: P=%b | Expected: P=%d",
                 673,
                 
                 P
                 , 
                 
                 2375
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110101; B = 7'b0001000; // Expected: {'P': 936}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110101; B = 7'b0001000; | Outputs: P=%b | Expected: P=%d",
                 674,
                 
                 P
                 , 
                 
                 936
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011001; B = 7'b0011000; // Expected: {'P': 2136}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011001; B = 7'b0011000; | Outputs: P=%b | Expected: P=%d",
                 675,
                 
                 P
                 , 
                 
                 2136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111111; B = 7'b0000011; // Expected: {'P': 189}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111111; B = 7'b0000011; | Outputs: P=%b | Expected: P=%d",
                 676,
                 
                 P
                 , 
                 
                 189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100011; B = 7'b1100111; // Expected: {'P': 10197}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100011; B = 7'b1100111; | Outputs: P=%b | Expected: P=%d",
                 677,
                 
                 P
                 , 
                 
                 10197
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110111; B = 7'b1110100; // Expected: {'P': 6380}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110111; B = 7'b1110100; | Outputs: P=%b | Expected: P=%d",
                 678,
                 
                 P
                 , 
                 
                 6380
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000111; B = 7'b0001000; // Expected: {'P': 568}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000111; B = 7'b0001000; | Outputs: P=%b | Expected: P=%d",
                 679,
                 
                 P
                 , 
                 
                 568
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101011; B = 7'b0101010; // Expected: {'P': 1806}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101011; B = 7'b0101010; | Outputs: P=%b | Expected: P=%d",
                 680,
                 
                 P
                 , 
                 
                 1806
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100110; B = 7'b1110110; // Expected: {'P': 4484}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100110; B = 7'b1110110; | Outputs: P=%b | Expected: P=%d",
                 681,
                 
                 P
                 , 
                 
                 4484
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110110; B = 7'b0010000; // Expected: {'P': 1888}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110110; B = 7'b0010000; | Outputs: P=%b | Expected: P=%d",
                 682,
                 
                 P
                 , 
                 
                 1888
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110110; B = 7'b0110010; // Expected: {'P': 2700}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110110; B = 7'b0110010; | Outputs: P=%b | Expected: P=%d",
                 683,
                 
                 P
                 , 
                 
                 2700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011100; B = 7'b1010101; // Expected: {'P': 2380}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011100; B = 7'b1010101; | Outputs: P=%b | Expected: P=%d",
                 684,
                 
                 P
                 , 
                 
                 2380
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001011; B = 7'b0101111; // Expected: {'P': 3525}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001011; B = 7'b0101111; | Outputs: P=%b | Expected: P=%d",
                 685,
                 
                 P
                 , 
                 
                 3525
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110111; B = 7'b1110100; // Expected: {'P': 13804}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110111; B = 7'b1110100; | Outputs: P=%b | Expected: P=%d",
                 686,
                 
                 P
                 , 
                 
                 13804
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100101; B = 7'b0000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100101; B = 7'b0000000; | Outputs: P=%b | Expected: P=%d",
                 687,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010010; B = 7'b0111000; // Expected: {'P': 4592}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010010; B = 7'b0111000; | Outputs: P=%b | Expected: P=%d",
                 688,
                 
                 P
                 , 
                 
                 4592
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111100; B = 7'b1000010; // Expected: {'P': 8184}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111100; B = 7'b1000010; | Outputs: P=%b | Expected: P=%d",
                 689,
                 
                 P
                 , 
                 
                 8184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101001; B = 7'b0001011; // Expected: {'P': 1155}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101001; B = 7'b0001011; | Outputs: P=%b | Expected: P=%d",
                 690,
                 
                 P
                 , 
                 
                 1155
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101110; B = 7'b1100000; // Expected: {'P': 10560}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101110; B = 7'b1100000; | Outputs: P=%b | Expected: P=%d",
                 691,
                 
                 P
                 , 
                 
                 10560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110010; B = 7'b0000011; // Expected: {'P': 150}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110010; B = 7'b0000011; | Outputs: P=%b | Expected: P=%d",
                 692,
                 
                 P
                 , 
                 
                 150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111101; B = 7'b0110001; // Expected: {'P': 2989}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111101; B = 7'b0110001; | Outputs: P=%b | Expected: P=%d",
                 693,
                 
                 P
                 , 
                 
                 2989
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010100; B = 7'b0000110; // Expected: {'P': 120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010100; B = 7'b0000110; | Outputs: P=%b | Expected: P=%d",
                 694,
                 
                 P
                 , 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011001; B = 7'b1110101; // Expected: {'P': 10413}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011001; B = 7'b1110101; | Outputs: P=%b | Expected: P=%d",
                 695,
                 
                 P
                 , 
                 
                 10413
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101110; B = 7'b0101110; // Expected: {'P': 5060}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101110; B = 7'b0101110; | Outputs: P=%b | Expected: P=%d",
                 696,
                 
                 P
                 , 
                 
                 5060
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010000; B = 7'b1100011; // Expected: {'P': 7920}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010000; B = 7'b1100011; | Outputs: P=%b | Expected: P=%d",
                 697,
                 
                 P
                 , 
                 
                 7920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101000; B = 7'b1110110; // Expected: {'P': 4720}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101000; B = 7'b1110110; | Outputs: P=%b | Expected: P=%d",
                 698,
                 
                 P
                 , 
                 
                 4720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011110; B = 7'b1000001; // Expected: {'P': 1950}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011110; B = 7'b1000001; | Outputs: P=%b | Expected: P=%d",
                 699,
                 
                 P
                 , 
                 
                 1950
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101110; B = 7'b0001111; // Expected: {'P': 690}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101110; B = 7'b0001111; | Outputs: P=%b | Expected: P=%d",
                 700,
                 
                 P
                 , 
                 
                 690
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100010; B = 7'b1101111; // Expected: {'P': 10878}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100010; B = 7'b1101111; | Outputs: P=%b | Expected: P=%d",
                 701,
                 
                 P
                 , 
                 
                 10878
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011011; B = 7'b1010110; // Expected: {'P': 7826}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011011; B = 7'b1010110; | Outputs: P=%b | Expected: P=%d",
                 702,
                 
                 P
                 , 
                 
                 7826
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100000; B = 7'b1111011; // Expected: {'P': 11808}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100000; B = 7'b1111011; | Outputs: P=%b | Expected: P=%d",
                 703,
                 
                 P
                 , 
                 
                 11808
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101101; B = 7'b0111001; // Expected: {'P': 6213}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101101; B = 7'b0111001; | Outputs: P=%b | Expected: P=%d",
                 704,
                 
                 P
                 , 
                 
                 6213
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111110; B = 7'b1110110; // Expected: {'P': 14868}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111110; B = 7'b1110110; | Outputs: P=%b | Expected: P=%d",
                 705,
                 
                 P
                 , 
                 
                 14868
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011010; B = 7'b0001100; // Expected: {'P': 1080}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011010; B = 7'b0001100; | Outputs: P=%b | Expected: P=%d",
                 706,
                 
                 P
                 , 
                 
                 1080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110010; B = 7'b1101111; // Expected: {'P': 12654}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110010; B = 7'b1101111; | Outputs: P=%b | Expected: P=%d",
                 707,
                 
                 P
                 , 
                 
                 12654
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010110; B = 7'b1001011; // Expected: {'P': 6450}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010110; B = 7'b1001011; | Outputs: P=%b | Expected: P=%d",
                 708,
                 
                 P
                 , 
                 
                 6450
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001011; B = 7'b0110010; // Expected: {'P': 550}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001011; B = 7'b0110010; | Outputs: P=%b | Expected: P=%d",
                 709,
                 
                 P
                 , 
                 
                 550
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101010; B = 7'b1001100; // Expected: {'P': 3192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101010; B = 7'b1001100; | Outputs: P=%b | Expected: P=%d",
                 710,
                 
                 P
                 , 
                 
                 3192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100100; B = 7'b0010111; // Expected: {'P': 2300}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100100; B = 7'b0010111; | Outputs: P=%b | Expected: P=%d",
                 711,
                 
                 P
                 , 
                 
                 2300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010011; B = 7'b0011010; // Expected: {'P': 2158}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010011; B = 7'b0011010; | Outputs: P=%b | Expected: P=%d",
                 712,
                 
                 P
                 , 
                 
                 2158
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000001; B = 7'b1101001; // Expected: {'P': 105}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000001; B = 7'b1101001; | Outputs: P=%b | Expected: P=%d",
                 713,
                 
                 P
                 , 
                 
                 105
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111001; B = 7'b0011101; // Expected: {'P': 3509}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111001; B = 7'b0011101; | Outputs: P=%b | Expected: P=%d",
                 714,
                 
                 P
                 , 
                 
                 3509
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101010; B = 7'b0010101; // Expected: {'P': 882}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101010; B = 7'b0010101; | Outputs: P=%b | Expected: P=%d",
                 715,
                 
                 P
                 , 
                 
                 882
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011011; B = 7'b0100001; // Expected: {'P': 3003}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011011; B = 7'b0100001; | Outputs: P=%b | Expected: P=%d",
                 716,
                 
                 P
                 , 
                 
                 3003
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110110; B = 7'b0110011; // Expected: {'P': 6018}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110110; B = 7'b0110011; | Outputs: P=%b | Expected: P=%d",
                 717,
                 
                 P
                 , 
                 
                 6018
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110000; B = 7'b1110111; // Expected: {'P': 5712}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110000; B = 7'b1110111; | Outputs: P=%b | Expected: P=%d",
                 718,
                 
                 P
                 , 
                 
                 5712
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100111; B = 7'b0100100; // Expected: {'P': 3708}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100111; B = 7'b0100100; | Outputs: P=%b | Expected: P=%d",
                 719,
                 
                 P
                 , 
                 
                 3708
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100011; B = 7'b1010111; // Expected: {'P': 3045}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100011; B = 7'b1010111; | Outputs: P=%b | Expected: P=%d",
                 720,
                 
                 P
                 , 
                 
                 3045
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110101; B = 7'b0101010; // Expected: {'P': 4914}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110101; B = 7'b0101010; | Outputs: P=%b | Expected: P=%d",
                 721,
                 
                 P
                 , 
                 
                 4914
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010010; B = 7'b1001011; // Expected: {'P': 1350}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010010; B = 7'b1001011; | Outputs: P=%b | Expected: P=%d",
                 722,
                 
                 P
                 , 
                 
                 1350
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111011; B = 7'b1001100; // Expected: {'P': 9348}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111011; B = 7'b1001100; | Outputs: P=%b | Expected: P=%d",
                 723,
                 
                 P
                 , 
                 
                 9348
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001010; B = 7'b1100111; // Expected: {'P': 1030}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001010; B = 7'b1100111; | Outputs: P=%b | Expected: P=%d",
                 724,
                 
                 P
                 , 
                 
                 1030
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111000; B = 7'b0000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111000; B = 7'b0000000; | Outputs: P=%b | Expected: P=%d",
                 725,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101100; B = 7'b1101011; // Expected: {'P': 11556}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101100; B = 7'b1101011; | Outputs: P=%b | Expected: P=%d",
                 726,
                 
                 P
                 , 
                 
                 11556
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111111; B = 7'b0101101; // Expected: {'P': 2835}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111111; B = 7'b0101101; | Outputs: P=%b | Expected: P=%d",
                 727,
                 
                 P
                 , 
                 
                 2835
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111100; B = 7'b1010000; // Expected: {'P': 9920}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111100; B = 7'b1010000; | Outputs: P=%b | Expected: P=%d",
                 728,
                 
                 P
                 , 
                 
                 9920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010110; B = 7'b0100001; // Expected: {'P': 2838}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010110; B = 7'b0100001; | Outputs: P=%b | Expected: P=%d",
                 729,
                 
                 P
                 , 
                 
                 2838
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111101; B = 7'b1110011; // Expected: {'P': 7015}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111101; B = 7'b1110011; | Outputs: P=%b | Expected: P=%d",
                 730,
                 
                 P
                 , 
                 
                 7015
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001000; B = 7'b0101000; // Expected: {'P': 320}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001000; B = 7'b0101000; | Outputs: P=%b | Expected: P=%d",
                 731,
                 
                 P
                 , 
                 
                 320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010110; B = 7'b1110110; // Expected: {'P': 10148}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010110; B = 7'b1110110; | Outputs: P=%b | Expected: P=%d",
                 732,
                 
                 P
                 , 
                 
                 10148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100110; B = 7'b0000110; // Expected: {'P': 228}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100110; B = 7'b0000110; | Outputs: P=%b | Expected: P=%d",
                 733,
                 
                 P
                 , 
                 
                 228
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011011; B = 7'b1001101; // Expected: {'P': 7007}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011011; B = 7'b1001101; | Outputs: P=%b | Expected: P=%d",
                 734,
                 
                 P
                 , 
                 
                 7007
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110000; B = 7'b0111000; // Expected: {'P': 6272}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110000; B = 7'b0111000; | Outputs: P=%b | Expected: P=%d",
                 735,
                 
                 P
                 , 
                 
                 6272
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101111; B = 7'b0100011; // Expected: {'P': 3885}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101111; B = 7'b0100011; | Outputs: P=%b | Expected: P=%d",
                 736,
                 
                 P
                 , 
                 
                 3885
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110011; B = 7'b0011100; // Expected: {'P': 3220}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110011; B = 7'b0011100; | Outputs: P=%b | Expected: P=%d",
                 737,
                 
                 P
                 , 
                 
                 3220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000100; B = 7'b1011100; // Expected: {'P': 368}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000100; B = 7'b1011100; | Outputs: P=%b | Expected: P=%d",
                 738,
                 
                 P
                 , 
                 
                 368
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001111; B = 7'b1111110; // Expected: {'P': 1890}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001111; B = 7'b1111110; | Outputs: P=%b | Expected: P=%d",
                 739,
                 
                 P
                 , 
                 
                 1890
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100101; B = 7'b1010111; // Expected: {'P': 3219}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100101; B = 7'b1010111; | Outputs: P=%b | Expected: P=%d",
                 740,
                 
                 P
                 , 
                 
                 3219
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100001; B = 7'b0101010; // Expected: {'P': 1386}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100001; B = 7'b0101010; | Outputs: P=%b | Expected: P=%d",
                 741,
                 
                 P
                 , 
                 
                 1386
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001111; B = 7'b1110011; // Expected: {'P': 1725}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001111; B = 7'b1110011; | Outputs: P=%b | Expected: P=%d",
                 742,
                 
                 P
                 , 
                 
                 1725
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101001; B = 7'b0100110; // Expected: {'P': 1558}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101001; B = 7'b0100110; | Outputs: P=%b | Expected: P=%d",
                 743,
                 
                 P
                 , 
                 
                 1558
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101100; B = 7'b0010101; // Expected: {'P': 2268}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101100; B = 7'b0010101; | Outputs: P=%b | Expected: P=%d",
                 744,
                 
                 P
                 , 
                 
                 2268
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101101; B = 7'b1100010; // Expected: {'P': 4410}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101101; B = 7'b1100010; | Outputs: P=%b | Expected: P=%d",
                 745,
                 
                 P
                 , 
                 
                 4410
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110101; B = 7'b0010111; // Expected: {'P': 2691}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110101; B = 7'b0010111; | Outputs: P=%b | Expected: P=%d",
                 746,
                 
                 P
                 , 
                 
                 2691
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000111; B = 7'b0010000; // Expected: {'P': 1136}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000111; B = 7'b0010000; | Outputs: P=%b | Expected: P=%d",
                 747,
                 
                 P
                 , 
                 
                 1136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010000; B = 7'b0001010; // Expected: {'P': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010000; B = 7'b0001010; | Outputs: P=%b | Expected: P=%d",
                 748,
                 
                 P
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101101; B = 7'b1110110; // Expected: {'P': 12862}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101101; B = 7'b1110110; | Outputs: P=%b | Expected: P=%d",
                 749,
                 
                 P
                 , 
                 
                 12862
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111011; B = 7'b1111100; // Expected: {'P': 7316}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111011; B = 7'b1111100; | Outputs: P=%b | Expected: P=%d",
                 750,
                 
                 P
                 , 
                 
                 7316
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100110; B = 7'b1010101; // Expected: {'P': 3230}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100110; B = 7'b1010101; | Outputs: P=%b | Expected: P=%d",
                 751,
                 
                 P
                 , 
                 
                 3230
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101110; B = 7'b0110101; // Expected: {'P': 2438}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101110; B = 7'b0110101; | Outputs: P=%b | Expected: P=%d",
                 752,
                 
                 P
                 , 
                 
                 2438
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000101; B = 7'b1110011; // Expected: {'P': 575}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000101; B = 7'b1110011; | Outputs: P=%b | Expected: P=%d",
                 753,
                 
                 P
                 , 
                 
                 575
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000100; B = 7'b1001101; // Expected: {'P': 308}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000100; B = 7'b1001101; | Outputs: P=%b | Expected: P=%d",
                 754,
                 
                 P
                 , 
                 
                 308
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111110; B = 7'b0000100; // Expected: {'P': 504}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111110; B = 7'b0000100; | Outputs: P=%b | Expected: P=%d",
                 755,
                 
                 P
                 , 
                 
                 504
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110110; B = 7'b0001111; // Expected: {'P': 810}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110110; B = 7'b0001111; | Outputs: P=%b | Expected: P=%d",
                 756,
                 
                 P
                 , 
                 
                 810
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100111; B = 7'b1000101; // Expected: {'P': 2691}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100111; B = 7'b1000101; | Outputs: P=%b | Expected: P=%d",
                 757,
                 
                 P
                 , 
                 
                 2691
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101101; B = 7'b0110000; // Expected: {'P': 5232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101101; B = 7'b0110000; | Outputs: P=%b | Expected: P=%d",
                 758,
                 
                 P
                 , 
                 
                 5232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101110; B = 7'b0011010; // Expected: {'P': 2860}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101110; B = 7'b0011010; | Outputs: P=%b | Expected: P=%d",
                 759,
                 
                 P
                 , 
                 
                 2860
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111111; B = 7'b1001101; // Expected: {'P': 4851}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111111; B = 7'b1001101; | Outputs: P=%b | Expected: P=%d",
                 760,
                 
                 P
                 , 
                 
                 4851
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111001; B = 7'b1110111; // Expected: {'P': 14399}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111001; B = 7'b1110111; | Outputs: P=%b | Expected: P=%d",
                 761,
                 
                 P
                 , 
                 
                 14399
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110101; B = 7'b1001110; // Expected: {'P': 4134}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110101; B = 7'b1001110; | Outputs: P=%b | Expected: P=%d",
                 762,
                 
                 P
                 , 
                 
                 4134
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010010; B = 7'b0000010; // Expected: {'P': 164}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010010; B = 7'b0000010; | Outputs: P=%b | Expected: P=%d",
                 763,
                 
                 P
                 , 
                 
                 164
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001100; B = 7'b1010110; // Expected: {'P': 6536}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001100; B = 7'b1010110; | Outputs: P=%b | Expected: P=%d",
                 764,
                 
                 P
                 , 
                 
                 6536
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100011; B = 7'b0000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100011; B = 7'b0000000; | Outputs: P=%b | Expected: P=%d",
                 765,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011001; B = 7'b1010100; // Expected: {'P': 2100}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011001; B = 7'b1010100; | Outputs: P=%b | Expected: P=%d",
                 766,
                 
                 P
                 , 
                 
                 2100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000001; B = 7'b1011011; // Expected: {'P': 5915}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000001; B = 7'b1011011; | Outputs: P=%b | Expected: P=%d",
                 767,
                 
                 P
                 , 
                 
                 5915
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101001; B = 7'b0010010; // Expected: {'P': 738}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101001; B = 7'b0010010; | Outputs: P=%b | Expected: P=%d",
                 768,
                 
                 P
                 , 
                 
                 738
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011010; B = 7'b0101010; // Expected: {'P': 3780}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011010; B = 7'b0101010; | Outputs: P=%b | Expected: P=%d",
                 769,
                 
                 P
                 , 
                 
                 3780
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110111; B = 7'b0001101; // Expected: {'P': 1547}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110111; B = 7'b0001101; | Outputs: P=%b | Expected: P=%d",
                 770,
                 
                 P
                 , 
                 
                 1547
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100011; B = 7'b0101111; // Expected: {'P': 1645}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100011; B = 7'b0101111; | Outputs: P=%b | Expected: P=%d",
                 771,
                 
                 P
                 , 
                 
                 1645
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000100; B = 7'b0000110; // Expected: {'P': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000100; B = 7'b0000110; | Outputs: P=%b | Expected: P=%d",
                 772,
                 
                 P
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101000; B = 7'b1000110; // Expected: {'P': 7280}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101000; B = 7'b1000110; | Outputs: P=%b | Expected: P=%d",
                 773,
                 
                 P
                 , 
                 
                 7280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111000; B = 7'b0111010; // Expected: {'P': 3248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111000; B = 7'b0111010; | Outputs: P=%b | Expected: P=%d",
                 774,
                 
                 P
                 , 
                 
                 3248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100110; B = 7'b1011010; // Expected: {'P': 3420}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100110; B = 7'b1011010; | Outputs: P=%b | Expected: P=%d",
                 775,
                 
                 P
                 , 
                 
                 3420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110001; B = 7'b0010011; // Expected: {'P': 931}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110001; B = 7'b0010011; | Outputs: P=%b | Expected: P=%d",
                 776,
                 
                 P
                 , 
                 
                 931
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111100; B = 7'b0001110; // Expected: {'P': 840}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111100; B = 7'b0001110; | Outputs: P=%b | Expected: P=%d",
                 777,
                 
                 P
                 , 
                 
                 840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110110; B = 7'b1000100; // Expected: {'P': 8024}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110110; B = 7'b1000100; | Outputs: P=%b | Expected: P=%d",
                 778,
                 
                 P
                 , 
                 
                 8024
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100001; B = 7'b1111010; // Expected: {'P': 11834}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100001; B = 7'b1111010; | Outputs: P=%b | Expected: P=%d",
                 779,
                 
                 P
                 , 
                 
                 11834
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110000; B = 7'b1011001; // Expected: {'P': 4272}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110000; B = 7'b1011001; | Outputs: P=%b | Expected: P=%d",
                 780,
                 
                 P
                 , 
                 
                 4272
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000000; B = 7'b1010001; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000000; B = 7'b1010001; | Outputs: P=%b | Expected: P=%d",
                 781,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100000; B = 7'b1011011; // Expected: {'P': 2912}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100000; B = 7'b1011011; | Outputs: P=%b | Expected: P=%d",
                 782,
                 
                 P
                 , 
                 
                 2912
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110110; B = 7'b1110111; // Expected: {'P': 14042}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110110; B = 7'b1110111; | Outputs: P=%b | Expected: P=%d",
                 783,
                 
                 P
                 , 
                 
                 14042
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100110; B = 7'b0001100; // Expected: {'P': 456}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100110; B = 7'b0001100; | Outputs: P=%b | Expected: P=%d",
                 784,
                 
                 P
                 , 
                 
                 456
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101000; B = 7'b1000010; // Expected: {'P': 2640}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101000; B = 7'b1000010; | Outputs: P=%b | Expected: P=%d",
                 785,
                 
                 P
                 , 
                 
                 2640
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110100; B = 7'b0011000; // Expected: {'P': 1248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110100; B = 7'b0011000; | Outputs: P=%b | Expected: P=%d",
                 786,
                 
                 P
                 , 
                 
                 1248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000001; B = 7'b0001011; // Expected: {'P': 715}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000001; B = 7'b0001011; | Outputs: P=%b | Expected: P=%d",
                 787,
                 
                 P
                 , 
                 
                 715
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111001; B = 7'b0101111; // Expected: {'P': 2679}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111001; B = 7'b0101111; | Outputs: P=%b | Expected: P=%d",
                 788,
                 
                 P
                 , 
                 
                 2679
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010010; B = 7'b0001111; // Expected: {'P': 270}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010010; B = 7'b0001111; | Outputs: P=%b | Expected: P=%d",
                 789,
                 
                 P
                 , 
                 
                 270
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101001; B = 7'b1110001; // Expected: {'P': 4633}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101001; B = 7'b1110001; | Outputs: P=%b | Expected: P=%d",
                 790,
                 
                 P
                 , 
                 
                 4633
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001000; B = 7'b0000001; // Expected: {'P': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001000; B = 7'b0000001; | Outputs: P=%b | Expected: P=%d",
                 791,
                 
                 P
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010100; B = 7'b0111001; // Expected: {'P': 1140}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010100; B = 7'b0111001; | Outputs: P=%b | Expected: P=%d",
                 792,
                 
                 P
                 , 
                 
                 1140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001101; B = 7'b1011000; // Expected: {'P': 1144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001101; B = 7'b1011000; | Outputs: P=%b | Expected: P=%d",
                 793,
                 
                 P
                 , 
                 
                 1144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101000; B = 7'b1110001; // Expected: {'P': 11752}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101000; B = 7'b1110001; | Outputs: P=%b | Expected: P=%d",
                 794,
                 
                 P
                 , 
                 
                 11752
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100110; B = 7'b1001001; // Expected: {'P': 7446}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100110; B = 7'b1001001; | Outputs: P=%b | Expected: P=%d",
                 795,
                 
                 P
                 , 
                 
                 7446
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101011; B = 7'b0110011; // Expected: {'P': 2193}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101011; B = 7'b0110011; | Outputs: P=%b | Expected: P=%d",
                 796,
                 
                 P
                 , 
                 
                 2193
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110110; B = 7'b0011100; // Expected: {'P': 3304}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110110; B = 7'b0011100; | Outputs: P=%b | Expected: P=%d",
                 797,
                 
                 P
                 , 
                 
                 3304
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101011; B = 7'b0110010; // Expected: {'P': 2150}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101011; B = 7'b0110010; | Outputs: P=%b | Expected: P=%d",
                 798,
                 
                 P
                 , 
                 
                 2150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111100; B = 7'b1110001; // Expected: {'P': 6780}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111100; B = 7'b1110001; | Outputs: P=%b | Expected: P=%d",
                 799,
                 
                 P
                 , 
                 
                 6780
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010101; B = 7'b0001011; // Expected: {'P': 935}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010101; B = 7'b0001011; | Outputs: P=%b | Expected: P=%d",
                 800,
                 
                 P
                 , 
                 
                 935
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001110; B = 7'b0110110; // Expected: {'P': 756}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001110; B = 7'b0110110; | Outputs: P=%b | Expected: P=%d",
                 801,
                 
                 P
                 , 
                 
                 756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010111; B = 7'b1101111; // Expected: {'P': 2553}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010111; B = 7'b1101111; | Outputs: P=%b | Expected: P=%d",
                 802,
                 
                 P
                 , 
                 
                 2553
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010010; B = 7'b0101010; // Expected: {'P': 3444}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010010; B = 7'b0101010; | Outputs: P=%b | Expected: P=%d",
                 803,
                 
                 P
                 , 
                 
                 3444
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100000; B = 7'b1110111; // Expected: {'P': 3808}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100000; B = 7'b1110111; | Outputs: P=%b | Expected: P=%d",
                 804,
                 
                 P
                 , 
                 
                 3808
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000010; B = 7'b0100011; // Expected: {'P': 2310}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000010; B = 7'b0100011; | Outputs: P=%b | Expected: P=%d",
                 805,
                 
                 P
                 , 
                 
                 2310
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000101; B = 7'b1111100; // Expected: {'P': 620}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000101; B = 7'b1111100; | Outputs: P=%b | Expected: P=%d",
                 806,
                 
                 P
                 , 
                 
                 620
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001111; B = 7'b1000111; // Expected: {'P': 5609}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001111; B = 7'b1000111; | Outputs: P=%b | Expected: P=%d",
                 807,
                 
                 P
                 , 
                 
                 5609
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111110; B = 7'b1110011; // Expected: {'P': 7130}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111110; B = 7'b1110011; | Outputs: P=%b | Expected: P=%d",
                 808,
                 
                 P
                 , 
                 
                 7130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110101; B = 7'b0011110; // Expected: {'P': 1590}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110101; B = 7'b0011110; | Outputs: P=%b | Expected: P=%d",
                 809,
                 
                 P
                 , 
                 
                 1590
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101110; B = 7'b0111101; // Expected: {'P': 6710}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101110; B = 7'b0111101; | Outputs: P=%b | Expected: P=%d",
                 810,
                 
                 P
                 , 
                 
                 6710
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101001; B = 7'b0101111; // Expected: {'P': 1927}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101001; B = 7'b0101111; | Outputs: P=%b | Expected: P=%d",
                 811,
                 
                 P
                 , 
                 
                 1927
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001110; B = 7'b1101001; // Expected: {'P': 1470}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001110; B = 7'b1101001; | Outputs: P=%b | Expected: P=%d",
                 812,
                 
                 P
                 , 
                 
                 1470
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101110; B = 7'b0001001; // Expected: {'P': 414}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101110; B = 7'b0001001; | Outputs: P=%b | Expected: P=%d",
                 813,
                 
                 P
                 , 
                 
                 414
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110010; B = 7'b0100001; // Expected: {'P': 1650}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110010; B = 7'b0100001; | Outputs: P=%b | Expected: P=%d",
                 814,
                 
                 P
                 , 
                 
                 1650
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011001; B = 7'b0111001; // Expected: {'P': 1425}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011001; B = 7'b0111001; | Outputs: P=%b | Expected: P=%d",
                 815,
                 
                 P
                 , 
                 
                 1425
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011001; B = 7'b1100101; // Expected: {'P': 2525}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011001; B = 7'b1100101; | Outputs: P=%b | Expected: P=%d",
                 816,
                 
                 P
                 , 
                 
                 2525
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100101; B = 7'b1000010; // Expected: {'P': 2442}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100101; B = 7'b1000010; | Outputs: P=%b | Expected: P=%d",
                 817,
                 
                 P
                 , 
                 
                 2442
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000011; B = 7'b0111100; // Expected: {'P': 180}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000011; B = 7'b0111100; | Outputs: P=%b | Expected: P=%d",
                 818,
                 
                 P
                 , 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001111; B = 7'b1101101; // Expected: {'P': 1635}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001111; B = 7'b1101101; | Outputs: P=%b | Expected: P=%d",
                 819,
                 
                 P
                 , 
                 
                 1635
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000001; B = 7'b0101011; // Expected: {'P': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000001; B = 7'b0101011; | Outputs: P=%b | Expected: P=%d",
                 820,
                 
                 P
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000001; B = 7'b0101101; // Expected: {'P': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000001; B = 7'b0101101; | Outputs: P=%b | Expected: P=%d",
                 821,
                 
                 P
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101110; B = 7'b0110111; // Expected: {'P': 2530}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101110; B = 7'b0110111; | Outputs: P=%b | Expected: P=%d",
                 822,
                 
                 P
                 , 
                 
                 2530
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010100; B = 7'b1110011; // Expected: {'P': 2300}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010100; B = 7'b1110011; | Outputs: P=%b | Expected: P=%d",
                 823,
                 
                 P
                 , 
                 
                 2300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000010; B = 7'b0100111; // Expected: {'P': 2574}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000010; B = 7'b0100111; | Outputs: P=%b | Expected: P=%d",
                 824,
                 
                 P
                 , 
                 
                 2574
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110010; B = 7'b0101101; // Expected: {'P': 5130}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110010; B = 7'b0101101; | Outputs: P=%b | Expected: P=%d",
                 825,
                 
                 P
                 , 
                 
                 5130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100001; B = 7'b0001110; // Expected: {'P': 1358}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100001; B = 7'b0001110; | Outputs: P=%b | Expected: P=%d",
                 826,
                 
                 P
                 , 
                 
                 1358
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011000; B = 7'b1111010; // Expected: {'P': 10736}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011000; B = 7'b1111010; | Outputs: P=%b | Expected: P=%d",
                 827,
                 
                 P
                 , 
                 
                 10736
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101100; B = 7'b0010100; // Expected: {'P': 2160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101100; B = 7'b0010100; | Outputs: P=%b | Expected: P=%d",
                 828,
                 
                 P
                 , 
                 
                 2160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000100; B = 7'b0111000; // Expected: {'P': 3808}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000100; B = 7'b0111000; | Outputs: P=%b | Expected: P=%d",
                 829,
                 
                 P
                 , 
                 
                 3808
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111000; B = 7'b1001100; // Expected: {'P': 9120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111000; B = 7'b1001100; | Outputs: P=%b | Expected: P=%d",
                 830,
                 
                 P
                 , 
                 
                 9120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110001; B = 7'b0010111; // Expected: {'P': 2599}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110001; B = 7'b0010111; | Outputs: P=%b | Expected: P=%d",
                 831,
                 
                 P
                 , 
                 
                 2599
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110101; B = 7'b0111100; // Expected: {'P': 7020}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110101; B = 7'b0111100; | Outputs: P=%b | Expected: P=%d",
                 832,
                 
                 P
                 , 
                 
                 7020
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000101; B = 7'b1001101; // Expected: {'P': 385}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000101; B = 7'b1001101; | Outputs: P=%b | Expected: P=%d",
                 833,
                 
                 P
                 , 
                 
                 385
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111101; B = 7'b1001100; // Expected: {'P': 9500}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111101; B = 7'b1001100; | Outputs: P=%b | Expected: P=%d",
                 834,
                 
                 P
                 , 
                 
                 9500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010011; B = 7'b1110110; // Expected: {'P': 2242}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010011; B = 7'b1110110; | Outputs: P=%b | Expected: P=%d",
                 835,
                 
                 P
                 , 
                 
                 2242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000110; B = 7'b0000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000110; B = 7'b0000000; | Outputs: P=%b | Expected: P=%d",
                 836,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101000; B = 7'b1100000; // Expected: {'P': 9984}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101000; B = 7'b1100000; | Outputs: P=%b | Expected: P=%d",
                 837,
                 
                 P
                 , 
                 
                 9984
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010010; B = 7'b0000001; // Expected: {'P': 82}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010010; B = 7'b0000001; | Outputs: P=%b | Expected: P=%d",
                 838,
                 
                 P
                 , 
                 
                 82
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100011; B = 7'b1000000; // Expected: {'P': 6336}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100011; B = 7'b1000000; | Outputs: P=%b | Expected: P=%d",
                 839,
                 
                 P
                 , 
                 
                 6336
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001101; B = 7'b1100000; // Expected: {'P': 7392}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001101; B = 7'b1100000; | Outputs: P=%b | Expected: P=%d",
                 840,
                 
                 P
                 , 
                 
                 7392
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110011; B = 7'b1011101; // Expected: {'P': 4743}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110011; B = 7'b1011101; | Outputs: P=%b | Expected: P=%d",
                 841,
                 
                 P
                 , 
                 
                 4743
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111011; B = 7'b0011001; // Expected: {'P': 3075}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111011; B = 7'b0011001; | Outputs: P=%b | Expected: P=%d",
                 842,
                 
                 P
                 , 
                 
                 3075
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110011; B = 7'b1100011; // Expected: {'P': 11385}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110011; B = 7'b1100011; | Outputs: P=%b | Expected: P=%d",
                 843,
                 
                 P
                 , 
                 
                 11385
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010100; B = 7'b1111110; // Expected: {'P': 2520}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010100; B = 7'b1111110; | Outputs: P=%b | Expected: P=%d",
                 844,
                 
                 P
                 , 
                 
                 2520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100100; B = 7'b1111100; // Expected: {'P': 12400}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100100; B = 7'b1111100; | Outputs: P=%b | Expected: P=%d",
                 845,
                 
                 P
                 , 
                 
                 12400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100110; B = 7'b1000110; // Expected: {'P': 7140}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100110; B = 7'b1000110; | Outputs: P=%b | Expected: P=%d",
                 846,
                 
                 P
                 , 
                 
                 7140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110111; B = 7'b0010111; // Expected: {'P': 2737}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110111; B = 7'b0010111; | Outputs: P=%b | Expected: P=%d",
                 847,
                 
                 P
                 , 
                 
                 2737
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001110; B = 7'b1111110; // Expected: {'P': 9828}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001110; B = 7'b1111110; | Outputs: P=%b | Expected: P=%d",
                 848,
                 
                 P
                 , 
                 
                 9828
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111110; B = 7'b1000100; // Expected: {'P': 4216}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111110; B = 7'b1000100; | Outputs: P=%b | Expected: P=%d",
                 849,
                 
                 P
                 , 
                 
                 4216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010000; B = 7'b1110101; // Expected: {'P': 9360}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010000; B = 7'b1110101; | Outputs: P=%b | Expected: P=%d",
                 850,
                 
                 P
                 , 
                 
                 9360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000000; B = 7'b1100000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000000; B = 7'b1100000; | Outputs: P=%b | Expected: P=%d",
                 851,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010111; B = 7'b0011110; // Expected: {'P': 690}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010111; B = 7'b0011110; | Outputs: P=%b | Expected: P=%d",
                 852,
                 
                 P
                 , 
                 
                 690
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111111; B = 7'b1110101; // Expected: {'P': 7371}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111111; B = 7'b1110101; | Outputs: P=%b | Expected: P=%d",
                 853,
                 
                 P
                 , 
                 
                 7371
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111110; B = 7'b1100100; // Expected: {'P': 12600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111110; B = 7'b1100100; | Outputs: P=%b | Expected: P=%d",
                 854,
                 
                 P
                 , 
                 
                 12600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001000; B = 7'b1111110; // Expected: {'P': 9072}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001000; B = 7'b1111110; | Outputs: P=%b | Expected: P=%d",
                 855,
                 
                 P
                 , 
                 
                 9072
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011111; B = 7'b0101001; // Expected: {'P': 3895}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011111; B = 7'b0101001; | Outputs: P=%b | Expected: P=%d",
                 856,
                 
                 P
                 , 
                 
                 3895
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100001; B = 7'b0101011; // Expected: {'P': 1419}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100001; B = 7'b0101011; | Outputs: P=%b | Expected: P=%d",
                 857,
                 
                 P
                 , 
                 
                 1419
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100010; B = 7'b1011011; // Expected: {'P': 8918}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100010; B = 7'b1011011; | Outputs: P=%b | Expected: P=%d",
                 858,
                 
                 P
                 , 
                 
                 8918
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001010; B = 7'b0111010; // Expected: {'P': 580}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001010; B = 7'b0111010; | Outputs: P=%b | Expected: P=%d",
                 859,
                 
                 P
                 , 
                 
                 580
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011001; B = 7'b0000101; // Expected: {'P': 445}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011001; B = 7'b0000101; | Outputs: P=%b | Expected: P=%d",
                 860,
                 
                 P
                 , 
                 
                 445
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101101; B = 7'b1010001; // Expected: {'P': 3645}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101101; B = 7'b1010001; | Outputs: P=%b | Expected: P=%d",
                 861,
                 
                 P
                 , 
                 
                 3645
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101010; B = 7'b0110110; // Expected: {'P': 2268}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101010; B = 7'b0110110; | Outputs: P=%b | Expected: P=%d",
                 862,
                 
                 P
                 , 
                 
                 2268
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100101; B = 7'b1010111; // Expected: {'P': 8787}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100101; B = 7'b1010111; | Outputs: P=%b | Expected: P=%d",
                 863,
                 
                 P
                 , 
                 
                 8787
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111101; B = 7'b0001000; // Expected: {'P': 1000}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111101; B = 7'b0001000; | Outputs: P=%b | Expected: P=%d",
                 864,
                 
                 P
                 , 
                 
                 1000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000010; B = 7'b1011000; // Expected: {'P': 176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000010; B = 7'b1011000; | Outputs: P=%b | Expected: P=%d",
                 865,
                 
                 P
                 , 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101101; B = 7'b0000010; // Expected: {'P': 218}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101101; B = 7'b0000010; | Outputs: P=%b | Expected: P=%d",
                 866,
                 
                 P
                 , 
                 
                 218
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011100; B = 7'b1100010; // Expected: {'P': 9016}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011100; B = 7'b1100010; | Outputs: P=%b | Expected: P=%d",
                 867,
                 
                 P
                 , 
                 
                 9016
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001100; B = 7'b1010111; // Expected: {'P': 6612}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001100; B = 7'b1010111; | Outputs: P=%b | Expected: P=%d",
                 868,
                 
                 P
                 , 
                 
                 6612
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011011; B = 7'b1111110; // Expected: {'P': 11466}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011011; B = 7'b1111110; | Outputs: P=%b | Expected: P=%d",
                 869,
                 
                 P
                 , 
                 
                 11466
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011011; B = 7'b0011111; // Expected: {'P': 837}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011011; B = 7'b0011111; | Outputs: P=%b | Expected: P=%d",
                 870,
                 
                 P
                 , 
                 
                 837
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000011; B = 7'b0010111; // Expected: {'P': 1541}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000011; B = 7'b0010111; | Outputs: P=%b | Expected: P=%d",
                 871,
                 
                 P
                 , 
                 
                 1541
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111110; B = 7'b0111011; // Expected: {'P': 7434}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111110; B = 7'b0111011; | Outputs: P=%b | Expected: P=%d",
                 872,
                 
                 P
                 , 
                 
                 7434
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101101; B = 7'b0011101; // Expected: {'P': 3161}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101101; B = 7'b0011101; | Outputs: P=%b | Expected: P=%d",
                 873,
                 
                 P
                 , 
                 
                 3161
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111001; B = 7'b0101010; // Expected: {'P': 5082}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111001; B = 7'b0101010; | Outputs: P=%b | Expected: P=%d",
                 874,
                 
                 P
                 , 
                 
                 5082
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000001; B = 7'b1100011; // Expected: {'P': 99}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000001; B = 7'b1100011; | Outputs: P=%b | Expected: P=%d",
                 875,
                 
                 P
                 , 
                 
                 99
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000001; B = 7'b1110000; // Expected: {'P': 112}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000001; B = 7'b1110000; | Outputs: P=%b | Expected: P=%d",
                 876,
                 
                 P
                 , 
                 
                 112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011001; B = 7'b0110111; // Expected: {'P': 1375}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011001; B = 7'b0110111; | Outputs: P=%b | Expected: P=%d",
                 877,
                 
                 P
                 , 
                 
                 1375
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000011; B = 7'b0000100; // Expected: {'P': 268}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000011; B = 7'b0000100; | Outputs: P=%b | Expected: P=%d",
                 878,
                 
                 P
                 , 
                 
                 268
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000010; B = 7'b0110110; // Expected: {'P': 108}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000010; B = 7'b0110110; | Outputs: P=%b | Expected: P=%d",
                 879,
                 
                 P
                 , 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100110; B = 7'b1001111; // Expected: {'P': 3002}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100110; B = 7'b1001111; | Outputs: P=%b | Expected: P=%d",
                 880,
                 
                 P
                 , 
                 
                 3002
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100111; B = 7'b0111001; // Expected: {'P': 5871}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100111; B = 7'b0111001; | Outputs: P=%b | Expected: P=%d",
                 881,
                 
                 P
                 , 
                 
                 5871
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111010; B = 7'b1111011; // Expected: {'P': 15006}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111010; B = 7'b1111011; | Outputs: P=%b | Expected: P=%d",
                 882,
                 
                 P
                 , 
                 
                 15006
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000010; B = 7'b1011001; // Expected: {'P': 5874}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000010; B = 7'b1011001; | Outputs: P=%b | Expected: P=%d",
                 883,
                 
                 P
                 , 
                 
                 5874
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011010; B = 7'b1011001; // Expected: {'P': 8010}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011010; B = 7'b1011001; | Outputs: P=%b | Expected: P=%d",
                 884,
                 
                 P
                 , 
                 
                 8010
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110100; B = 7'b0111011; // Expected: {'P': 3068}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110100; B = 7'b0111011; | Outputs: P=%b | Expected: P=%d",
                 885,
                 
                 P
                 , 
                 
                 3068
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011001; B = 7'b1110000; // Expected: {'P': 9968}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011001; B = 7'b1110000; | Outputs: P=%b | Expected: P=%d",
                 886,
                 
                 P
                 , 
                 
                 9968
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010101; B = 7'b0100101; // Expected: {'P': 777}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010101; B = 7'b0100101; | Outputs: P=%b | Expected: P=%d",
                 887,
                 
                 P
                 , 
                 
                 777
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001000; B = 7'b1110100; // Expected: {'P': 8352}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001000; B = 7'b1110100; | Outputs: P=%b | Expected: P=%d",
                 888,
                 
                 P
                 , 
                 
                 8352
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100111; B = 7'b0011100; // Expected: {'P': 1092}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100111; B = 7'b0011100; | Outputs: P=%b | Expected: P=%d",
                 889,
                 
                 P
                 , 
                 
                 1092
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001000; B = 7'b1100111; // Expected: {'P': 7416}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001000; B = 7'b1100111; | Outputs: P=%b | Expected: P=%d",
                 890,
                 
                 P
                 , 
                 
                 7416
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101000; B = 7'b1111010; // Expected: {'P': 4880}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101000; B = 7'b1111010; | Outputs: P=%b | Expected: P=%d",
                 891,
                 
                 P
                 , 
                 
                 4880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111001; B = 7'b0011101; // Expected: {'P': 1653}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111001; B = 7'b0011101; | Outputs: P=%b | Expected: P=%d",
                 892,
                 
                 P
                 , 
                 
                 1653
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010010; B = 7'b1101111; // Expected: {'P': 1998}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010010; B = 7'b1101111; | Outputs: P=%b | Expected: P=%d",
                 893,
                 
                 P
                 , 
                 
                 1998
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010000; B = 7'b0110010; // Expected: {'P': 4000}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010000; B = 7'b0110010; | Outputs: P=%b | Expected: P=%d",
                 894,
                 
                 P
                 , 
                 
                 4000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000001; B = 7'b0011111; // Expected: {'P': 31}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000001; B = 7'b0011111; | Outputs: P=%b | Expected: P=%d",
                 895,
                 
                 P
                 , 
                 
                 31
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101100; B = 7'b0010110; // Expected: {'P': 2376}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101100; B = 7'b0010110; | Outputs: P=%b | Expected: P=%d",
                 896,
                 
                 P
                 , 
                 
                 2376
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111011; B = 7'b0011100; // Expected: {'P': 3444}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111011; B = 7'b0011100; | Outputs: P=%b | Expected: P=%d",
                 897,
                 
                 P
                 , 
                 
                 3444
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100110; B = 7'b1001000; // Expected: {'P': 2736}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100110; B = 7'b1001000; | Outputs: P=%b | Expected: P=%d",
                 898,
                 
                 P
                 , 
                 
                 2736
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010001; B = 7'b0000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010001; B = 7'b0000000; | Outputs: P=%b | Expected: P=%d",
                 899,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010100; B = 7'b1111110; // Expected: {'P': 10584}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010100; B = 7'b1111110; | Outputs: P=%b | Expected: P=%d",
                 900,
                 
                 P
                 , 
                 
                 10584
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011010; B = 7'b1001101; // Expected: {'P': 2002}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011010; B = 7'b1001101; | Outputs: P=%b | Expected: P=%d",
                 901,
                 
                 P
                 , 
                 
                 2002
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001110; B = 7'b1011110; // Expected: {'P': 7332}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001110; B = 7'b1011110; | Outputs: P=%b | Expected: P=%d",
                 902,
                 
                 P
                 , 
                 
                 7332
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100111; B = 7'b1101001; // Expected: {'P': 4095}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100111; B = 7'b1101001; | Outputs: P=%b | Expected: P=%d",
                 903,
                 
                 P
                 , 
                 
                 4095
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100011; B = 7'b0100100; // Expected: {'P': 3564}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100011; B = 7'b0100100; | Outputs: P=%b | Expected: P=%d",
                 904,
                 
                 P
                 , 
                 
                 3564
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111010; B = 7'b1110100; // Expected: {'P': 14152}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111010; B = 7'b1110100; | Outputs: P=%b | Expected: P=%d",
                 905,
                 
                 P
                 , 
                 
                 14152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110010; B = 7'b1010100; // Expected: {'P': 4200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110010; B = 7'b1010100; | Outputs: P=%b | Expected: P=%d",
                 906,
                 
                 P
                 , 
                 
                 4200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010011; B = 7'b0110110; // Expected: {'P': 1026}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010011; B = 7'b0110110; | Outputs: P=%b | Expected: P=%d",
                 907,
                 
                 P
                 , 
                 
                 1026
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001110; B = 7'b0100110; // Expected: {'P': 532}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001110; B = 7'b0100110; | Outputs: P=%b | Expected: P=%d",
                 908,
                 
                 P
                 , 
                 
                 532
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011110; B = 7'b1111000; // Expected: {'P': 11280}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011110; B = 7'b1111000; | Outputs: P=%b | Expected: P=%d",
                 909,
                 
                 P
                 , 
                 
                 11280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010101; B = 7'b1110010; // Expected: {'P': 2394}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010101; B = 7'b1110010; | Outputs: P=%b | Expected: P=%d",
                 910,
                 
                 P
                 , 
                 
                 2394
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001101; B = 7'b0100110; // Expected: {'P': 2926}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001101; B = 7'b0100110; | Outputs: P=%b | Expected: P=%d",
                 911,
                 
                 P
                 , 
                 
                 2926
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110000; B = 7'b1101000; // Expected: {'P': 11648}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110000; B = 7'b1101000; | Outputs: P=%b | Expected: P=%d",
                 912,
                 
                 P
                 , 
                 
                 11648
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001001; B = 7'b1010000; // Expected: {'P': 5840}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001001; B = 7'b1010000; | Outputs: P=%b | Expected: P=%d",
                 913,
                 
                 P
                 , 
                 
                 5840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110111; B = 7'b1100100; // Expected: {'P': 5500}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110111; B = 7'b1100100; | Outputs: P=%b | Expected: P=%d",
                 914,
                 
                 P
                 , 
                 
                 5500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110100; B = 7'b0011011; // Expected: {'P': 1404}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110100; B = 7'b0011011; | Outputs: P=%b | Expected: P=%d",
                 915,
                 
                 P
                 , 
                 
                 1404
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011001; B = 7'b0010100; // Expected: {'P': 500}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011001; B = 7'b0010100; | Outputs: P=%b | Expected: P=%d",
                 916,
                 
                 P
                 , 
                 
                 500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100110; B = 7'b1100100; // Expected: {'P': 10200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100110; B = 7'b1100100; | Outputs: P=%b | Expected: P=%d",
                 917,
                 
                 P
                 , 
                 
                 10200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010001; B = 7'b0011011; // Expected: {'P': 2187}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010001; B = 7'b0011011; | Outputs: P=%b | Expected: P=%d",
                 918,
                 
                 P
                 , 
                 
                 2187
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010000; B = 7'b1000100; // Expected: {'P': 5440}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010000; B = 7'b1000100; | Outputs: P=%b | Expected: P=%d",
                 919,
                 
                 P
                 , 
                 
                 5440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111101; B = 7'b1001000; // Expected: {'P': 9000}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111101; B = 7'b1001000; | Outputs: P=%b | Expected: P=%d",
                 920,
                 
                 P
                 , 
                 
                 9000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001100; B = 7'b0110111; // Expected: {'P': 660}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001100; B = 7'b0110111; | Outputs: P=%b | Expected: P=%d",
                 921,
                 
                 P
                 , 
                 
                 660
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111000; B = 7'b1010100; // Expected: {'P': 4704}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111000; B = 7'b1010100; | Outputs: P=%b | Expected: P=%d",
                 922,
                 
                 P
                 , 
                 
                 4704
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110100; B = 7'b0010111; // Expected: {'P': 2668}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110100; B = 7'b0010111; | Outputs: P=%b | Expected: P=%d",
                 923,
                 
                 P
                 , 
                 
                 2668
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101011; B = 7'b0010010; // Expected: {'P': 774}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101011; B = 7'b0010010; | Outputs: P=%b | Expected: P=%d",
                 924,
                 
                 P
                 , 
                 
                 774
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010011; B = 7'b0110111; // Expected: {'P': 4565}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010011; B = 7'b0110111; | Outputs: P=%b | Expected: P=%d",
                 925,
                 
                 P
                 , 
                 
                 4565
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011001; B = 7'b0011001; // Expected: {'P': 2225}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011001; B = 7'b0011001; | Outputs: P=%b | Expected: P=%d",
                 926,
                 
                 P
                 , 
                 
                 2225
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110000; B = 7'b0101010; // Expected: {'P': 2016}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110000; B = 7'b0101010; | Outputs: P=%b | Expected: P=%d",
                 927,
                 
                 P
                 , 
                 
                 2016
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010101; B = 7'b0001000; // Expected: {'P': 168}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010101; B = 7'b0001000; | Outputs: P=%b | Expected: P=%d",
                 928,
                 
                 P
                 , 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001001; B = 7'b1100001; // Expected: {'P': 7081}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001001; B = 7'b1100001; | Outputs: P=%b | Expected: P=%d",
                 929,
                 
                 P
                 , 
                 
                 7081
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110100; B = 7'b0111010; // Expected: {'P': 3016}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110100; B = 7'b0111010; | Outputs: P=%b | Expected: P=%d",
                 930,
                 
                 P
                 , 
                 
                 3016
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110111; B = 7'b1101110; // Expected: {'P': 6050}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110111; B = 7'b1101110; | Outputs: P=%b | Expected: P=%d",
                 931,
                 
                 P
                 , 
                 
                 6050
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110100; B = 7'b1111101; // Expected: {'P': 14500}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110100; B = 7'b1111101; | Outputs: P=%b | Expected: P=%d",
                 932,
                 
                 P
                 , 
                 
                 14500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000011; B = 7'b1010000; // Expected: {'P': 5360}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000011; B = 7'b1010000; | Outputs: P=%b | Expected: P=%d",
                 933,
                 
                 P
                 , 
                 
                 5360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000010; B = 7'b1111000; // Expected: {'P': 7920}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000010; B = 7'b1111000; | Outputs: P=%b | Expected: P=%d",
                 934,
                 
                 P
                 , 
                 
                 7920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000010; B = 7'b1011110; // Expected: {'P': 188}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000010; B = 7'b1011110; | Outputs: P=%b | Expected: P=%d",
                 935,
                 
                 P
                 , 
                 
                 188
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101100; B = 7'b0110101; // Expected: {'P': 5724}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101100; B = 7'b0110101; | Outputs: P=%b | Expected: P=%d",
                 936,
                 
                 P
                 , 
                 
                 5724
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010100; B = 7'b0100110; // Expected: {'P': 3192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010100; B = 7'b0100110; | Outputs: P=%b | Expected: P=%d",
                 937,
                 
                 P
                 , 
                 
                 3192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111100; B = 7'b0001001; // Expected: {'P': 540}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111100; B = 7'b0001001; | Outputs: P=%b | Expected: P=%d",
                 938,
                 
                 P
                 , 
                 
                 540
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011011; B = 7'b1101001; // Expected: {'P': 2835}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011011; B = 7'b1101001; | Outputs: P=%b | Expected: P=%d",
                 939,
                 
                 P
                 , 
                 
                 2835
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101010; B = 7'b1111100; // Expected: {'P': 13144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101010; B = 7'b1111100; | Outputs: P=%b | Expected: P=%d",
                 940,
                 
                 P
                 , 
                 
                 13144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010101; B = 7'b0111010; // Expected: {'P': 4930}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010101; B = 7'b0111010; | Outputs: P=%b | Expected: P=%d",
                 941,
                 
                 P
                 , 
                 
                 4930
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100010; B = 7'b1101101; // Expected: {'P': 10682}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100010; B = 7'b1101101; | Outputs: P=%b | Expected: P=%d",
                 942,
                 
                 P
                 , 
                 
                 10682
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110110; B = 7'b1010000; // Expected: {'P': 9440}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110110; B = 7'b1010000; | Outputs: P=%b | Expected: P=%d",
                 943,
                 
                 P
                 , 
                 
                 9440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111111; B = 7'b1110101; // Expected: {'P': 14859}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111111; B = 7'b1110101; | Outputs: P=%b | Expected: P=%d",
                 944,
                 
                 P
                 , 
                 
                 14859
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011101; B = 7'b0011110; // Expected: {'P': 2790}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011101; B = 7'b0011110; | Outputs: P=%b | Expected: P=%d",
                 945,
                 
                 P
                 , 
                 
                 2790
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110111; B = 7'b0100100; // Expected: {'P': 1980}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110111; B = 7'b0100100; | Outputs: P=%b | Expected: P=%d",
                 946,
                 
                 P
                 , 
                 
                 1980
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000110; B = 7'b0101010; // Expected: {'P': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000110; B = 7'b0101010; | Outputs: P=%b | Expected: P=%d",
                 947,
                 
                 P
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100110; B = 7'b0111111; // Expected: {'P': 2394}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100110; B = 7'b0111111; | Outputs: P=%b | Expected: P=%d",
                 948,
                 
                 P
                 , 
                 
                 2394
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111111; B = 7'b1011111; // Expected: {'P': 12065}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111111; B = 7'b1011111; | Outputs: P=%b | Expected: P=%d",
                 949,
                 
                 P
                 , 
                 
                 12065
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011101; B = 7'b0101101; // Expected: {'P': 4185}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011101; B = 7'b0101101; | Outputs: P=%b | Expected: P=%d",
                 950,
                 
                 P
                 , 
                 
                 4185
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101100; B = 7'b1011100; // Expected: {'P': 4048}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101100; B = 7'b1011100; | Outputs: P=%b | Expected: P=%d",
                 951,
                 
                 P
                 , 
                 
                 4048
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001110; B = 7'b0011001; // Expected: {'P': 350}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001110; B = 7'b0011001; | Outputs: P=%b | Expected: P=%d",
                 952,
                 
                 P
                 , 
                 
                 350
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000000; B = 7'b1100000; // Expected: {'P': 6144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000000; B = 7'b1100000; | Outputs: P=%b | Expected: P=%d",
                 953,
                 
                 P
                 , 
                 
                 6144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111011; B = 7'b1011000; // Expected: {'P': 10824}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111011; B = 7'b1011000; | Outputs: P=%b | Expected: P=%d",
                 954,
                 
                 P
                 , 
                 
                 10824
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110010; B = 7'b1101000; // Expected: {'P': 5200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110010; B = 7'b1101000; | Outputs: P=%b | Expected: P=%d",
                 955,
                 
                 P
                 , 
                 
                 5200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001111; B = 7'b1001010; // Expected: {'P': 5846}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001111; B = 7'b1001010; | Outputs: P=%b | Expected: P=%d",
                 956,
                 
                 P
                 , 
                 
                 5846
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010000; B = 7'b1010001; // Expected: {'P': 6480}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010000; B = 7'b1010001; | Outputs: P=%b | Expected: P=%d",
                 957,
                 
                 P
                 , 
                 
                 6480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101010; B = 7'b0111101; // Expected: {'P': 6466}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101010; B = 7'b0111101; | Outputs: P=%b | Expected: P=%d",
                 958,
                 
                 P
                 , 
                 
                 6466
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100010; B = 7'b1101100; // Expected: {'P': 3672}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100010; B = 7'b1101100; | Outputs: P=%b | Expected: P=%d",
                 959,
                 
                 P
                 , 
                 
                 3672
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111101; B = 7'b1101110; // Expected: {'P': 6710}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111101; B = 7'b1101110; | Outputs: P=%b | Expected: P=%d",
                 960,
                 
                 P
                 , 
                 
                 6710
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110110; B = 7'b1000011; // Expected: {'P': 3618}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110110; B = 7'b1000011; | Outputs: P=%b | Expected: P=%d",
                 961,
                 
                 P
                 , 
                 
                 3618
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010001; B = 7'b0100010; // Expected: {'P': 2754}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010001; B = 7'b0100010; | Outputs: P=%b | Expected: P=%d",
                 962,
                 
                 P
                 , 
                 
                 2754
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101111; B = 7'b1110100; // Expected: {'P': 5452}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101111; B = 7'b1110100; | Outputs: P=%b | Expected: P=%d",
                 963,
                 
                 P
                 , 
                 
                 5452
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011010; B = 7'b0101101; // Expected: {'P': 1170}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011010; B = 7'b0101101; | Outputs: P=%b | Expected: P=%d",
                 964,
                 
                 P
                 , 
                 
                 1170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111100; B = 7'b1101011; // Expected: {'P': 13268}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111100; B = 7'b1101011; | Outputs: P=%b | Expected: P=%d",
                 965,
                 
                 P
                 , 
                 
                 13268
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111011; B = 7'b1000101; // Expected: {'P': 8487}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111011; B = 7'b1000101; | Outputs: P=%b | Expected: P=%d",
                 966,
                 
                 P
                 , 
                 
                 8487
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110100; B = 7'b0010100; // Expected: {'P': 1040}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110100; B = 7'b0010100; | Outputs: P=%b | Expected: P=%d",
                 967,
                 
                 P
                 , 
                 
                 1040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000001; B = 7'b0100100; // Expected: {'P': 36}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000001; B = 7'b0100100; | Outputs: P=%b | Expected: P=%d",
                 968,
                 
                 P
                 , 
                 
                 36
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001111; B = 7'b0100000; // Expected: {'P': 2528}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001111; B = 7'b0100000; | Outputs: P=%b | Expected: P=%d",
                 969,
                 
                 P
                 , 
                 
                 2528
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010001; B = 7'b0100100; // Expected: {'P': 612}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010001; B = 7'b0100100; | Outputs: P=%b | Expected: P=%d",
                 970,
                 
                 P
                 , 
                 
                 612
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010110; B = 7'b0010111; // Expected: {'P': 1978}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010110; B = 7'b0010111; | Outputs: P=%b | Expected: P=%d",
                 971,
                 
                 P
                 , 
                 
                 1978
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110010; B = 7'b1111100; // Expected: {'P': 14136}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110010; B = 7'b1111100; | Outputs: P=%b | Expected: P=%d",
                 972,
                 
                 P
                 , 
                 
                 14136
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110100; B = 7'b0111111; // Expected: {'P': 3276}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110100; B = 7'b0111111; | Outputs: P=%b | Expected: P=%d",
                 973,
                 
                 P
                 , 
                 
                 3276
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000111; B = 7'b1010010; // Expected: {'P': 574}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000111; B = 7'b1010010; | Outputs: P=%b | Expected: P=%d",
                 974,
                 
                 P
                 , 
                 
                 574
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111111; B = 7'b1001001; // Expected: {'P': 9271}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111111; B = 7'b1001001; | Outputs: P=%b | Expected: P=%d",
                 975,
                 
                 P
                 , 
                 
                 9271
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001010; B = 7'b1011000; // Expected: {'P': 6512}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001010; B = 7'b1011000; | Outputs: P=%b | Expected: P=%d",
                 976,
                 
                 P
                 , 
                 
                 6512
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011001; B = 7'b0000110; // Expected: {'P': 534}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011001; B = 7'b0000110; | Outputs: P=%b | Expected: P=%d",
                 977,
                 
                 P
                 , 
                 
                 534
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111010; B = 7'b1111000; // Expected: {'P': 6960}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111010; B = 7'b1111000; | Outputs: P=%b | Expected: P=%d",
                 978,
                 
                 P
                 , 
                 
                 6960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101110; B = 7'b0001101; // Expected: {'P': 598}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101110; B = 7'b0001101; | Outputs: P=%b | Expected: P=%d",
                 979,
                 
                 P
                 , 
                 
                 598
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000101; B = 7'b0010110; // Expected: {'P': 110}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000101; B = 7'b0010110; | Outputs: P=%b | Expected: P=%d",
                 980,
                 
                 P
                 , 
                 
                 110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101001; B = 7'b1001010; // Expected: {'P': 3034}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101001; B = 7'b1001010; | Outputs: P=%b | Expected: P=%d",
                 981,
                 
                 P
                 , 
                 
                 3034
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110011; B = 7'b0101110; // Expected: {'P': 2346}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110011; B = 7'b0101110; | Outputs: P=%b | Expected: P=%d",
                 982,
                 
                 P
                 , 
                 
                 2346
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011010; B = 7'b0011010; // Expected: {'P': 676}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011010; B = 7'b0011010; | Outputs: P=%b | Expected: P=%d",
                 983,
                 
                 P
                 , 
                 
                 676
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101011; B = 7'b1101000; // Expected: {'P': 11128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101011; B = 7'b1101000; | Outputs: P=%b | Expected: P=%d",
                 984,
                 
                 P
                 , 
                 
                 11128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010010; B = 7'b0110010; // Expected: {'P': 900}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010010; B = 7'b0110010; | Outputs: P=%b | Expected: P=%d",
                 985,
                 
                 P
                 , 
                 
                 900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110110; B = 7'b1000000; // Expected: {'P': 7552}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110110; B = 7'b1000000; | Outputs: P=%b | Expected: P=%d",
                 986,
                 
                 P
                 , 
                 
                 7552
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001011; B = 7'b1010000; // Expected: {'P': 6000}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001011; B = 7'b1010000; | Outputs: P=%b | Expected: P=%d",
                 987,
                 
                 P
                 , 
                 
                 6000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110101; B = 7'b0000001; // Expected: {'P': 117}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110101; B = 7'b0000001; | Outputs: P=%b | Expected: P=%d",
                 988,
                 
                 P
                 , 
                 
                 117
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101001; B = 7'b1000011; // Expected: {'P': 2747}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101001; B = 7'b1000011; | Outputs: P=%b | Expected: P=%d",
                 989,
                 
                 P
                 , 
                 
                 2747
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010010; B = 7'b0101001; // Expected: {'P': 738}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010010; B = 7'b0101001; | Outputs: P=%b | Expected: P=%d",
                 990,
                 
                 P
                 , 
                 
                 738
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100111; B = 7'b1101111; // Expected: {'P': 11433}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100111; B = 7'b1101111; | Outputs: P=%b | Expected: P=%d",
                 991,
                 
                 P
                 , 
                 
                 11433
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111111; B = 7'b0010100; // Expected: {'P': 1260}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111111; B = 7'b0010100; | Outputs: P=%b | Expected: P=%d",
                 992,
                 
                 P
                 , 
                 
                 1260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010001; B = 7'b1100100; // Expected: {'P': 1700}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010001; B = 7'b1100100; | Outputs: P=%b | Expected: P=%d",
                 993,
                 
                 P
                 , 
                 
                 1700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101001; B = 7'b0011100; // Expected: {'P': 1148}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101001; B = 7'b0011100; | Outputs: P=%b | Expected: P=%d",
                 994,
                 
                 P
                 , 
                 
                 1148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011001; B = 7'b0001101; // Expected: {'P': 1157}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011001; B = 7'b0001101; | Outputs: P=%b | Expected: P=%d",
                 995,
                 
                 P
                 , 
                 
                 1157
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110111; B = 7'b1110111; // Expected: {'P': 6545}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110111; B = 7'b1110111; | Outputs: P=%b | Expected: P=%d",
                 996,
                 
                 P
                 , 
                 
                 6545
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111101; B = 7'b1110000; // Expected: {'P': 6832}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111101; B = 7'b1110000; | Outputs: P=%b | Expected: P=%d",
                 997,
                 
                 P
                 , 
                 
                 6832
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001100; B = 7'b1001101; // Expected: {'P': 5852}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001100; B = 7'b1001101; | Outputs: P=%b | Expected: P=%d",
                 998,
                 
                 P
                 , 
                 
                 5852
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011100; B = 7'b1101010; // Expected: {'P': 9752}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011100; B = 7'b1101010; | Outputs: P=%b | Expected: P=%d",
                 999,
                 
                 P
                 , 
                 
                 9752
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011110; B = 7'b1001110; // Expected: {'P': 7332}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011110; B = 7'b1001110; | Outputs: P=%b | Expected: P=%d",
                 1000,
                 
                 P
                 , 
                 
                 7332
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001011; B = 7'b0101010; // Expected: {'P': 3150}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001011; B = 7'b0101010; | Outputs: P=%b | Expected: P=%d",
                 1001,
                 
                 P
                 , 
                 
                 3150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100010; B = 7'b0010001; // Expected: {'P': 578}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100010; B = 7'b0010001; | Outputs: P=%b | Expected: P=%d",
                 1002,
                 
                 P
                 , 
                 
                 578
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000110; B = 7'b0001110; // Expected: {'P': 980}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000110; B = 7'b0001110; | Outputs: P=%b | Expected: P=%d",
                 1003,
                 
                 P
                 , 
                 
                 980
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110110; B = 7'b0100001; // Expected: {'P': 3894}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110110; B = 7'b0100001; | Outputs: P=%b | Expected: P=%d",
                 1004,
                 
                 P
                 , 
                 
                 3894
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010111; B = 7'b1001000; // Expected: {'P': 6264}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010111; B = 7'b1001000; | Outputs: P=%b | Expected: P=%d",
                 1005,
                 
                 P
                 , 
                 
                 6264
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101010; B = 7'b0110001; // Expected: {'P': 5194}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101010; B = 7'b0110001; | Outputs: P=%b | Expected: P=%d",
                 1006,
                 
                 P
                 , 
                 
                 5194
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110100; B = 7'b1101100; // Expected: {'P': 5616}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110100; B = 7'b1101100; | Outputs: P=%b | Expected: P=%d",
                 1007,
                 
                 P
                 , 
                 
                 5616
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101001; B = 7'b0000100; // Expected: {'P': 420}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101001; B = 7'b0000100; | Outputs: P=%b | Expected: P=%d",
                 1008,
                 
                 P
                 , 
                 
                 420
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111100; B = 7'b0100100; // Expected: {'P': 4464}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111100; B = 7'b0100100; | Outputs: P=%b | Expected: P=%d",
                 1009,
                 
                 P
                 , 
                 
                 4464
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000100; B = 7'b1011011; // Expected: {'P': 364}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000100; B = 7'b1011011; | Outputs: P=%b | Expected: P=%d",
                 1010,
                 
                 P
                 , 
                 
                 364
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111000; B = 7'b0000110; // Expected: {'P': 336}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111000; B = 7'b0000110; | Outputs: P=%b | Expected: P=%d",
                 1011,
                 
                 P
                 , 
                 
                 336
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000011; B = 7'b1111101; // Expected: {'P': 375}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000011; B = 7'b1111101; | Outputs: P=%b | Expected: P=%d",
                 1012,
                 
                 P
                 , 
                 
                 375
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111001; B = 7'b0010100; // Expected: {'P': 1140}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111001; B = 7'b0010100; | Outputs: P=%b | Expected: P=%d",
                 1013,
                 
                 P
                 , 
                 
                 1140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000011; B = 7'b1000011; // Expected: {'P': 4489}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000011; B = 7'b1000011; | Outputs: P=%b | Expected: P=%d",
                 1014,
                 
                 P
                 , 
                 
                 4489
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010110; B = 7'b1111111; // Expected: {'P': 2794}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010110; B = 7'b1111111; | Outputs: P=%b | Expected: P=%d",
                 1015,
                 
                 P
                 , 
                 
                 2794
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001111; B = 7'b1001111; // Expected: {'P': 6241}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001111; B = 7'b1001111; | Outputs: P=%b | Expected: P=%d",
                 1016,
                 
                 P
                 , 
                 
                 6241
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011111; B = 7'b1000000; // Expected: {'P': 6080}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011111; B = 7'b1000000; | Outputs: P=%b | Expected: P=%d",
                 1017,
                 
                 P
                 , 
                 
                 6080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100011; B = 7'b1101111; // Expected: {'P': 3885}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100011; B = 7'b1101111; | Outputs: P=%b | Expected: P=%d",
                 1018,
                 
                 P
                 , 
                 
                 3885
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010101; B = 7'b1101011; // Expected: {'P': 2247}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010101; B = 7'b1101011; | Outputs: P=%b | Expected: P=%d",
                 1019,
                 
                 P
                 , 
                 
                 2247
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111101; B = 7'b1111110; // Expected: {'P': 15750}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111101; B = 7'b1111110; | Outputs: P=%b | Expected: P=%d",
                 1020,
                 
                 P
                 , 
                 
                 15750
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010011; B = 7'b1111100; // Expected: {'P': 2356}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010011; B = 7'b1111100; | Outputs: P=%b | Expected: P=%d",
                 1021,
                 
                 P
                 , 
                 
                 2356
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100101; B = 7'b1100101; // Expected: {'P': 10201}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100101; B = 7'b1100101; | Outputs: P=%b | Expected: P=%d",
                 1022,
                 
                 P
                 , 
                 
                 10201
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110010; B = 7'b0110100; // Expected: {'P': 2600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110010; B = 7'b0110100; | Outputs: P=%b | Expected: P=%d",
                 1023,
                 
                 P
                 , 
                 
                 2600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110101; B = 7'b1100111; // Expected: {'P': 12051}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110101; B = 7'b1100111; | Outputs: P=%b | Expected: P=%d",
                 1024,
                 
                 P
                 , 
                 
                 12051
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000110; B = 7'b0100111; // Expected: {'P': 2730}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000110; B = 7'b0100111; | Outputs: P=%b | Expected: P=%d",
                 1025,
                 
                 P
                 , 
                 
                 2730
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101001; B = 7'b1011000; // Expected: {'P': 3608}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101001; B = 7'b1011000; | Outputs: P=%b | Expected: P=%d",
                 1026,
                 
                 P
                 , 
                 
                 3608
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010111; B = 7'b1011001; // Expected: {'P': 7743}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010111; B = 7'b1011001; | Outputs: P=%b | Expected: P=%d",
                 1027,
                 
                 P
                 , 
                 
                 7743
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100101; B = 7'b0111010; // Expected: {'P': 5858}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100101; B = 7'b0111010; | Outputs: P=%b | Expected: P=%d",
                 1028,
                 
                 P
                 , 
                 
                 5858
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100101; B = 7'b1100010; // Expected: {'P': 9898}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100101; B = 7'b1100010; | Outputs: P=%b | Expected: P=%d",
                 1029,
                 
                 P
                 , 
                 
                 9898
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001101; B = 7'b0000101; // Expected: {'P': 385}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001101; B = 7'b0000101; | Outputs: P=%b | Expected: P=%d",
                 1030,
                 
                 P
                 , 
                 
                 385
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011001; B = 7'b0111010; // Expected: {'P': 5162}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011001; B = 7'b0111010; | Outputs: P=%b | Expected: P=%d",
                 1031,
                 
                 P
                 , 
                 
                 5162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110010; B = 7'b0000110; // Expected: {'P': 684}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110010; B = 7'b0000110; | Outputs: P=%b | Expected: P=%d",
                 1032,
                 
                 P
                 , 
                 
                 684
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001001; B = 7'b1101010; // Expected: {'P': 954}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001001; B = 7'b1101010; | Outputs: P=%b | Expected: P=%d",
                 1033,
                 
                 P
                 , 
                 
                 954
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110010; B = 7'b0001100; // Expected: {'P': 600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110010; B = 7'b0001100; | Outputs: P=%b | Expected: P=%d",
                 1034,
                 
                 P
                 , 
                 
                 600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000101; B = 7'b1110000; // Expected: {'P': 560}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000101; B = 7'b1110000; | Outputs: P=%b | Expected: P=%d",
                 1035,
                 
                 P
                 , 
                 
                 560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010111; B = 7'b1001110; // Expected: {'P': 6786}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010111; B = 7'b1001110; | Outputs: P=%b | Expected: P=%d",
                 1036,
                 
                 P
                 , 
                 
                 6786
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000000; B = 7'b1011101; // Expected: {'P': 5952}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000000; B = 7'b1011101; | Outputs: P=%b | Expected: P=%d",
                 1037,
                 
                 P
                 , 
                 
                 5952
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110000; B = 7'b1101101; // Expected: {'P': 5232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110000; B = 7'b1101101; | Outputs: P=%b | Expected: P=%d",
                 1038,
                 
                 P
                 , 
                 
                 5232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110110; B = 7'b1001010; // Expected: {'P': 8732}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110110; B = 7'b1001010; | Outputs: P=%b | Expected: P=%d",
                 1039,
                 
                 P
                 , 
                 
                 8732
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000001; B = 7'b1010111; // Expected: {'P': 5655}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000001; B = 7'b1010111; | Outputs: P=%b | Expected: P=%d",
                 1040,
                 
                 P
                 , 
                 
                 5655
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010000; B = 7'b0001100; // Expected: {'P': 192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010000; B = 7'b0001100; | Outputs: P=%b | Expected: P=%d",
                 1041,
                 
                 P
                 , 
                 
                 192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100010; B = 7'b1100110; // Expected: {'P': 3468}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100010; B = 7'b1100110; | Outputs: P=%b | Expected: P=%d",
                 1042,
                 
                 P
                 , 
                 
                 3468
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100000; B = 7'b1101101; // Expected: {'P': 10464}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100000; B = 7'b1101101; | Outputs: P=%b | Expected: P=%d",
                 1043,
                 
                 P
                 , 
                 
                 10464
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000010; B = 7'b0101001; // Expected: {'P': 82}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000010; B = 7'b0101001; | Outputs: P=%b | Expected: P=%d",
                 1044,
                 
                 P
                 , 
                 
                 82
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010010; B = 7'b0000011; // Expected: {'P': 54}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010010; B = 7'b0000011; | Outputs: P=%b | Expected: P=%d",
                 1045,
                 
                 P
                 , 
                 
                 54
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100101; B = 7'b0001001; // Expected: {'P': 909}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100101; B = 7'b0001001; | Outputs: P=%b | Expected: P=%d",
                 1046,
                 
                 P
                 , 
                 
                 909
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010100; B = 7'b0101100; // Expected: {'P': 880}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010100; B = 7'b0101100; | Outputs: P=%b | Expected: P=%d",
                 1047,
                 
                 P
                 , 
                 
                 880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100011; B = 7'b0100100; // Expected: {'P': 1260}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100011; B = 7'b0100100; | Outputs: P=%b | Expected: P=%d",
                 1048,
                 
                 P
                 , 
                 
                 1260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110110; B = 7'b0111000; // Expected: {'P': 6608}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110110; B = 7'b0111000; | Outputs: P=%b | Expected: P=%d",
                 1049,
                 
                 P
                 , 
                 
                 6608
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001110; B = 7'b0001011; // Expected: {'P': 154}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001110; B = 7'b0001011; | Outputs: P=%b | Expected: P=%d",
                 1050,
                 
                 P
                 , 
                 
                 154
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001001; B = 7'b0010011; // Expected: {'P': 171}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001001; B = 7'b0010011; | Outputs: P=%b | Expected: P=%d",
                 1051,
                 
                 P
                 , 
                 
                 171
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111000; B = 7'b1101111; // Expected: {'P': 13320}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111000; B = 7'b1101111; | Outputs: P=%b | Expected: P=%d",
                 1052,
                 
                 P
                 , 
                 
                 13320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111010; B = 7'b1110000; // Expected: {'P': 6496}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111010; B = 7'b1110000; | Outputs: P=%b | Expected: P=%d",
                 1053,
                 
                 P
                 , 
                 
                 6496
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111100; B = 7'b1001110; // Expected: {'P': 9672}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111100; B = 7'b1001110; | Outputs: P=%b | Expected: P=%d",
                 1054,
                 
                 P
                 , 
                 
                 9672
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110011; B = 7'b1110111; // Expected: {'P': 13685}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110011; B = 7'b1110111; | Outputs: P=%b | Expected: P=%d",
                 1055,
                 
                 P
                 , 
                 
                 13685
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111010; B = 7'b1001100; // Expected: {'P': 4408}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111010; B = 7'b1001100; | Outputs: P=%b | Expected: P=%d",
                 1056,
                 
                 P
                 , 
                 
                 4408
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100110; B = 7'b0100101; // Expected: {'P': 1406}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100110; B = 7'b0100101; | Outputs: P=%b | Expected: P=%d",
                 1057,
                 
                 P
                 , 
                 
                 1406
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101000; B = 7'b0010000; // Expected: {'P': 640}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101000; B = 7'b0010000; | Outputs: P=%b | Expected: P=%d",
                 1058,
                 
                 P
                 , 
                 
                 640
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101110; B = 7'b0110110; // Expected: {'P': 2484}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101110; B = 7'b0110110; | Outputs: P=%b | Expected: P=%d",
                 1059,
                 
                 P
                 , 
                 
                 2484
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010011; B = 7'b1001101; // Expected: {'P': 1463}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010011; B = 7'b1001101; | Outputs: P=%b | Expected: P=%d",
                 1060,
                 
                 P
                 , 
                 
                 1463
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111110; B = 7'b1001011; // Expected: {'P': 4650}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111110; B = 7'b1001011; | Outputs: P=%b | Expected: P=%d",
                 1061,
                 
                 P
                 , 
                 
                 4650
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100000; B = 7'b0011101; // Expected: {'P': 2784}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100000; B = 7'b0011101; | Outputs: P=%b | Expected: P=%d",
                 1062,
                 
                 P
                 , 
                 
                 2784
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001101; B = 7'b0100111; // Expected: {'P': 3003}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001101; B = 7'b0100111; | Outputs: P=%b | Expected: P=%d",
                 1063,
                 
                 P
                 , 
                 
                 3003
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100000; B = 7'b0100110; // Expected: {'P': 3648}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100000; B = 7'b0100110; | Outputs: P=%b | Expected: P=%d",
                 1064,
                 
                 P
                 , 
                 
                 3648
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100010; B = 7'b0011000; // Expected: {'P': 816}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100010; B = 7'b0011000; | Outputs: P=%b | Expected: P=%d",
                 1065,
                 
                 P
                 , 
                 
                 816
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110000; B = 7'b0111100; // Expected: {'P': 2880}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110000; B = 7'b0111100; | Outputs: P=%b | Expected: P=%d",
                 1066,
                 
                 P
                 , 
                 
                 2880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011000; B = 7'b0000111; // Expected: {'P': 616}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011000; B = 7'b0000111; | Outputs: P=%b | Expected: P=%d",
                 1067,
                 
                 P
                 , 
                 
                 616
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111111; B = 7'b1011010; // Expected: {'P': 5670}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111111; B = 7'b1011010; | Outputs: P=%b | Expected: P=%d",
                 1068,
                 
                 P
                 , 
                 
                 5670
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111111; B = 7'b1110111; // Expected: {'P': 15113}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111111; B = 7'b1110111; | Outputs: P=%b | Expected: P=%d",
                 1069,
                 
                 P
                 , 
                 
                 15113
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100001; B = 7'b0100001; // Expected: {'P': 3201}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100001; B = 7'b0100001; | Outputs: P=%b | Expected: P=%d",
                 1070,
                 
                 P
                 , 
                 
                 3201
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011000; B = 7'b0100011; // Expected: {'P': 3080}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011000; B = 7'b0100011; | Outputs: P=%b | Expected: P=%d",
                 1071,
                 
                 P
                 , 
                 
                 3080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000000; B = 7'b1001010; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000000; B = 7'b1001010; | Outputs: P=%b | Expected: P=%d",
                 1072,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010011; B = 7'b0010110; // Expected: {'P': 418}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010011; B = 7'b0010110; | Outputs: P=%b | Expected: P=%d",
                 1073,
                 
                 P
                 , 
                 
                 418
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100111; B = 7'b0110010; // Expected: {'P': 1950}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100111; B = 7'b0110010; | Outputs: P=%b | Expected: P=%d",
                 1074,
                 
                 P
                 , 
                 
                 1950
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101001; B = 7'b1010101; // Expected: {'P': 8925}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101001; B = 7'b1010101; | Outputs: P=%b | Expected: P=%d",
                 1075,
                 
                 P
                 , 
                 
                 8925
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101101; B = 7'b0100111; // Expected: {'P': 1755}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101101; B = 7'b0100111; | Outputs: P=%b | Expected: P=%d",
                 1076,
                 
                 P
                 , 
                 
                 1755
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101110; B = 7'b1101110; // Expected: {'P': 5060}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101110; B = 7'b1101110; | Outputs: P=%b | Expected: P=%d",
                 1077,
                 
                 P
                 , 
                 
                 5060
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111011; B = 7'b1100010; // Expected: {'P': 12054}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111011; B = 7'b1100010; | Outputs: P=%b | Expected: P=%d",
                 1078,
                 
                 P
                 , 
                 
                 12054
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001101; B = 7'b0111010; // Expected: {'P': 754}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001101; B = 7'b0111010; | Outputs: P=%b | Expected: P=%d",
                 1079,
                 
                 P
                 , 
                 
                 754
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000110; B = 7'b0000111; // Expected: {'P': 490}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000110; B = 7'b0000111; | Outputs: P=%b | Expected: P=%d",
                 1080,
                 
                 P
                 , 
                 
                 490
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101100; B = 7'b1001101; // Expected: {'P': 8316}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101100; B = 7'b1001101; | Outputs: P=%b | Expected: P=%d",
                 1081,
                 
                 P
                 , 
                 
                 8316
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000110; B = 7'b0101110; // Expected: {'P': 3220}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000110; B = 7'b0101110; | Outputs: P=%b | Expected: P=%d",
                 1082,
                 
                 P
                 , 
                 
                 3220
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011101; B = 7'b0100010; // Expected: {'P': 3162}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011101; B = 7'b0100010; | Outputs: P=%b | Expected: P=%d",
                 1083,
                 
                 P
                 , 
                 
                 3162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101011; B = 7'b0001110; // Expected: {'P': 1498}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101011; B = 7'b0001110; | Outputs: P=%b | Expected: P=%d",
                 1084,
                 
                 P
                 , 
                 
                 1498
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110010; B = 7'b1001101; // Expected: {'P': 3850}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110010; B = 7'b1001101; | Outputs: P=%b | Expected: P=%d",
                 1085,
                 
                 P
                 , 
                 
                 3850
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000110; B = 7'b0000100; // Expected: {'P': 24}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000110; B = 7'b0000100; | Outputs: P=%b | Expected: P=%d",
                 1086,
                 
                 P
                 , 
                 
                 24
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001010; B = 7'b1001110; // Expected: {'P': 5772}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001010; B = 7'b1001110; | Outputs: P=%b | Expected: P=%d",
                 1087,
                 
                 P
                 , 
                 
                 5772
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110100; B = 7'b1011011; // Expected: {'P': 10556}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110100; B = 7'b1011011; | Outputs: P=%b | Expected: P=%d",
                 1088,
                 
                 P
                 , 
                 
                 10556
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110001; B = 7'b1000001; // Expected: {'P': 7345}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110001; B = 7'b1000001; | Outputs: P=%b | Expected: P=%d",
                 1089,
                 
                 P
                 , 
                 
                 7345
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111101; B = 7'b1110110; // Expected: {'P': 14750}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111101; B = 7'b1110110; | Outputs: P=%b | Expected: P=%d",
                 1090,
                 
                 P
                 , 
                 
                 14750
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010000; B = 7'b0101001; // Expected: {'P': 3280}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010000; B = 7'b0101001; | Outputs: P=%b | Expected: P=%d",
                 1091,
                 
                 P
                 , 
                 
                 3280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111100; B = 7'b1010001; // Expected: {'P': 4860}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111100; B = 7'b1010001; | Outputs: P=%b | Expected: P=%d",
                 1092,
                 
                 P
                 , 
                 
                 4860
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101100; B = 7'b1000110; // Expected: {'P': 7560}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101100; B = 7'b1000110; | Outputs: P=%b | Expected: P=%d",
                 1093,
                 
                 P
                 , 
                 
                 7560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010101; B = 7'b0001100; // Expected: {'P': 1020}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010101; B = 7'b0001100; | Outputs: P=%b | Expected: P=%d",
                 1094,
                 
                 P
                 , 
                 
                 1020
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001011; B = 7'b0101000; // Expected: {'P': 3000}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001011; B = 7'b0101000; | Outputs: P=%b | Expected: P=%d",
                 1095,
                 
                 P
                 , 
                 
                 3000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011101; B = 7'b0101011; // Expected: {'P': 3999}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011101; B = 7'b0101011; | Outputs: P=%b | Expected: P=%d",
                 1096,
                 
                 P
                 , 
                 
                 3999
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011100; B = 7'b0011101; // Expected: {'P': 812}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011100; B = 7'b0011101; | Outputs: P=%b | Expected: P=%d",
                 1097,
                 
                 P
                 , 
                 
                 812
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010101; B = 7'b1000011; // Expected: {'P': 1407}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010101; B = 7'b1000011; | Outputs: P=%b | Expected: P=%d",
                 1098,
                 
                 P
                 , 
                 
                 1407
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000111; B = 7'b1111010; // Expected: {'P': 8662}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000111; B = 7'b1111010; | Outputs: P=%b | Expected: P=%d",
                 1099,
                 
                 P
                 , 
                 
                 8662
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010011; B = 7'b1000111; // Expected: {'P': 5893}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010011; B = 7'b1000111; | Outputs: P=%b | Expected: P=%d",
                 1100,
                 
                 P
                 , 
                 
                 5893
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000110; B = 7'b0100010; // Expected: {'P': 204}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000110; B = 7'b0100010; | Outputs: P=%b | Expected: P=%d",
                 1101,
                 
                 P
                 , 
                 
                 204
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111101; B = 7'b0010100; // Expected: {'P': 2500}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111101; B = 7'b0010100; | Outputs: P=%b | Expected: P=%d",
                 1102,
                 
                 P
                 , 
                 
                 2500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100011; B = 7'b1011101; // Expected: {'P': 3255}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100011; B = 7'b1011101; | Outputs: P=%b | Expected: P=%d",
                 1103,
                 
                 P
                 , 
                 
                 3255
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110100; B = 7'b0011011; // Expected: {'P': 3132}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110100; B = 7'b0011011; | Outputs: P=%b | Expected: P=%d",
                 1104,
                 
                 P
                 , 
                 
                 3132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100101; B = 7'b0110011; // Expected: {'P': 5151}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100101; B = 7'b0110011; | Outputs: P=%b | Expected: P=%d",
                 1105,
                 
                 P
                 , 
                 
                 5151
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110010; B = 7'b0101100; // Expected: {'P': 2200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110010; B = 7'b0101100; | Outputs: P=%b | Expected: P=%d",
                 1106,
                 
                 P
                 , 
                 
                 2200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111001; B = 7'b1010001; // Expected: {'P': 4617}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111001; B = 7'b1010001; | Outputs: P=%b | Expected: P=%d",
                 1107,
                 
                 P
                 , 
                 
                 4617
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100000; B = 7'b1101110; // Expected: {'P': 10560}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100000; B = 7'b1101110; | Outputs: P=%b | Expected: P=%d",
                 1108,
                 
                 P
                 , 
                 
                 10560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101100; B = 7'b0001101; // Expected: {'P': 1404}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101100; B = 7'b0001101; | Outputs: P=%b | Expected: P=%d",
                 1109,
                 
                 P
                 , 
                 
                 1404
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100011; B = 7'b1100110; // Expected: {'P': 3570}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100011; B = 7'b1100110; | Outputs: P=%b | Expected: P=%d",
                 1110,
                 
                 P
                 , 
                 
                 3570
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100110; B = 7'b0101011; // Expected: {'P': 1634}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100110; B = 7'b0101011; | Outputs: P=%b | Expected: P=%d",
                 1111,
                 
                 P
                 , 
                 
                 1634
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110001; B = 7'b1110010; // Expected: {'P': 5586}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110001; B = 7'b1110010; | Outputs: P=%b | Expected: P=%d",
                 1112,
                 
                 P
                 , 
                 
                 5586
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101011; B = 7'b1000000; // Expected: {'P': 6848}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101011; B = 7'b1000000; | Outputs: P=%b | Expected: P=%d",
                 1113,
                 
                 P
                 , 
                 
                 6848
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101110; B = 7'b1010011; // Expected: {'P': 9130}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101110; B = 7'b1010011; | Outputs: P=%b | Expected: P=%d",
                 1114,
                 
                 P
                 , 
                 
                 9130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011000; B = 7'b0011000; // Expected: {'P': 2112}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011000; B = 7'b0011000; | Outputs: P=%b | Expected: P=%d",
                 1115,
                 
                 P
                 , 
                 
                 2112
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101111; B = 7'b1001010; // Expected: {'P': 3478}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101111; B = 7'b1001010; | Outputs: P=%b | Expected: P=%d",
                 1116,
                 
                 P
                 , 
                 
                 3478
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000101; B = 7'b0001100; // Expected: {'P': 60}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000101; B = 7'b0001100; | Outputs: P=%b | Expected: P=%d",
                 1117,
                 
                 P
                 , 
                 
                 60
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010001; B = 7'b1011100; // Expected: {'P': 1564}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010001; B = 7'b1011100; | Outputs: P=%b | Expected: P=%d",
                 1118,
                 
                 P
                 , 
                 
                 1564
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111101; B = 7'b0011111; // Expected: {'P': 1891}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111101; B = 7'b0011111; | Outputs: P=%b | Expected: P=%d",
                 1119,
                 
                 P
                 , 
                 
                 1891
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000010; B = 7'b0101100; // Expected: {'P': 88}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000010; B = 7'b0101100; | Outputs: P=%b | Expected: P=%d",
                 1120,
                 
                 P
                 , 
                 
                 88
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001010; B = 7'b0100110; // Expected: {'P': 2812}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001010; B = 7'b0100110; | Outputs: P=%b | Expected: P=%d",
                 1121,
                 
                 P
                 , 
                 
                 2812
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011000; B = 7'b1011100; // Expected: {'P': 8096}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011000; B = 7'b1011100; | Outputs: P=%b | Expected: P=%d",
                 1122,
                 
                 P
                 , 
                 
                 8096
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010011; B = 7'b1111101; // Expected: {'P': 2375}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010011; B = 7'b1111101; | Outputs: P=%b | Expected: P=%d",
                 1123,
                 
                 P
                 , 
                 
                 2375
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101011; B = 7'b0010000; // Expected: {'P': 1712}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101011; B = 7'b0010000; | Outputs: P=%b | Expected: P=%d",
                 1124,
                 
                 P
                 , 
                 
                 1712
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010001; B = 7'b0110001; // Expected: {'P': 833}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010001; B = 7'b0110001; | Outputs: P=%b | Expected: P=%d",
                 1125,
                 
                 P
                 , 
                 
                 833
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111111; B = 7'b0111100; // Expected: {'P': 7620}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111111; B = 7'b0111100; | Outputs: P=%b | Expected: P=%d",
                 1126,
                 
                 P
                 , 
                 
                 7620
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011010; B = 7'b0001010; // Expected: {'P': 260}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011010; B = 7'b0001010; | Outputs: P=%b | Expected: P=%d",
                 1127,
                 
                 P
                 , 
                 
                 260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011011; B = 7'b1010101; // Expected: {'P': 2295}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011011; B = 7'b1010101; | Outputs: P=%b | Expected: P=%d",
                 1128,
                 
                 P
                 , 
                 
                 2295
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111001; B = 7'b1011100; // Expected: {'P': 11132}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111001; B = 7'b1011100; | Outputs: P=%b | Expected: P=%d",
                 1129,
                 
                 P
                 , 
                 
                 11132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100000; B = 7'b0001010; // Expected: {'P': 320}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100000; B = 7'b0001010; | Outputs: P=%b | Expected: P=%d",
                 1130,
                 
                 P
                 , 
                 
                 320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110111; B = 7'b0011010; // Expected: {'P': 3094}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110111; B = 7'b0011010; | Outputs: P=%b | Expected: P=%d",
                 1131,
                 
                 P
                 , 
                 
                 3094
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111001; B = 7'b1010110; // Expected: {'P': 10406}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111001; B = 7'b1010110; | Outputs: P=%b | Expected: P=%d",
                 1132,
                 
                 P
                 , 
                 
                 10406
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100000; B = 7'b0010010; // Expected: {'P': 576}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100000; B = 7'b0010010; | Outputs: P=%b | Expected: P=%d",
                 1133,
                 
                 P
                 , 
                 
                 576
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011101; B = 7'b1010010; // Expected: {'P': 7626}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011101; B = 7'b1010010; | Outputs: P=%b | Expected: P=%d",
                 1134,
                 
                 P
                 , 
                 
                 7626
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111101; B = 7'b0010101; // Expected: {'P': 1281}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111101; B = 7'b0010101; | Outputs: P=%b | Expected: P=%d",
                 1135,
                 
                 P
                 , 
                 
                 1281
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011110; B = 7'b1101010; // Expected: {'P': 3180}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011110; B = 7'b1101010; | Outputs: P=%b | Expected: P=%d",
                 1136,
                 
                 P
                 , 
                 
                 3180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101110; B = 7'b1001101; // Expected: {'P': 8470}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101110; B = 7'b1001101; | Outputs: P=%b | Expected: P=%d",
                 1137,
                 
                 P
                 , 
                 
                 8470
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101100; B = 7'b1011010; // Expected: {'P': 9720}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101100; B = 7'b1011010; | Outputs: P=%b | Expected: P=%d",
                 1138,
                 
                 P
                 , 
                 
                 9720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111101; B = 7'b1101101; // Expected: {'P': 13625}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111101; B = 7'b1101101; | Outputs: P=%b | Expected: P=%d",
                 1139,
                 
                 P
                 , 
                 
                 13625
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111111; B = 7'b1110001; // Expected: {'P': 14351}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111111; B = 7'b1110001; | Outputs: P=%b | Expected: P=%d",
                 1140,
                 
                 P
                 , 
                 
                 14351
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100000; B = 7'b1110101; // Expected: {'P': 11232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100000; B = 7'b1110101; | Outputs: P=%b | Expected: P=%d",
                 1141,
                 
                 P
                 , 
                 
                 11232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110010; B = 7'b0011000; // Expected: {'P': 2736}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110010; B = 7'b0011000; | Outputs: P=%b | Expected: P=%d",
                 1142,
                 
                 P
                 , 
                 
                 2736
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100011; B = 7'b1011001; // Expected: {'P': 3115}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100011; B = 7'b1011001; | Outputs: P=%b | Expected: P=%d",
                 1143,
                 
                 P
                 , 
                 
                 3115
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111001; B = 7'b1111011; // Expected: {'P': 7011}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111001; B = 7'b1111011; | Outputs: P=%b | Expected: P=%d",
                 1144,
                 
                 P
                 , 
                 
                 7011
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011010; B = 7'b0010111; // Expected: {'P': 2070}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011010; B = 7'b0010111; | Outputs: P=%b | Expected: P=%d",
                 1145,
                 
                 P
                 , 
                 
                 2070
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010000; B = 7'b0101100; // Expected: {'P': 3520}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010000; B = 7'b0101100; | Outputs: P=%b | Expected: P=%d",
                 1146,
                 
                 P
                 , 
                 
                 3520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010010; B = 7'b0001100; // Expected: {'P': 984}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010010; B = 7'b0001100; | Outputs: P=%b | Expected: P=%d",
                 1147,
                 
                 P
                 , 
                 
                 984
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101000; B = 7'b1110110; // Expected: {'P': 12272}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101000; B = 7'b1110110; | Outputs: P=%b | Expected: P=%d",
                 1148,
                 
                 P
                 , 
                 
                 12272
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000101; B = 7'b1000111; // Expected: {'P': 355}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000101; B = 7'b1000111; | Outputs: P=%b | Expected: P=%d",
                 1149,
                 
                 P
                 , 
                 
                 355
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110110; B = 7'b1101101; // Expected: {'P': 12862}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110110; B = 7'b1101101; | Outputs: P=%b | Expected: P=%d",
                 1150,
                 
                 P
                 , 
                 
                 12862
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010011; B = 7'b1010101; // Expected: {'P': 7055}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010011; B = 7'b1010101; | Outputs: P=%b | Expected: P=%d",
                 1151,
                 
                 P
                 , 
                 
                 7055
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101011; B = 7'b1010001; // Expected: {'P': 3483}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101011; B = 7'b1010001; | Outputs: P=%b | Expected: P=%d",
                 1152,
                 
                 P
                 , 
                 
                 3483
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110001; B = 7'b1110100; // Expected: {'P': 13108}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110001; B = 7'b1110100; | Outputs: P=%b | Expected: P=%d",
                 1153,
                 
                 P
                 , 
                 
                 13108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000111; B = 7'b1111000; // Expected: {'P': 840}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000111; B = 7'b1111000; | Outputs: P=%b | Expected: P=%d",
                 1154,
                 
                 P
                 , 
                 
                 840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001101; B = 7'b1010100; // Expected: {'P': 1092}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001101; B = 7'b1010100; | Outputs: P=%b | Expected: P=%d",
                 1155,
                 
                 P
                 , 
                 
                 1092
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100111; B = 7'b1000010; // Expected: {'P': 2574}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100111; B = 7'b1000010; | Outputs: P=%b | Expected: P=%d",
                 1156,
                 
                 P
                 , 
                 
                 2574
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010110; B = 7'b0110101; // Expected: {'P': 1166}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010110; B = 7'b0110101; | Outputs: P=%b | Expected: P=%d",
                 1157,
                 
                 P
                 , 
                 
                 1166
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100010; B = 7'b0110001; // Expected: {'P': 1666}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100010; B = 7'b0110001; | Outputs: P=%b | Expected: P=%d",
                 1158,
                 
                 P
                 , 
                 
                 1666
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011101; B = 7'b0110001; // Expected: {'P': 4557}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011101; B = 7'b0110001; | Outputs: P=%b | Expected: P=%d",
                 1159,
                 
                 P
                 , 
                 
                 4557
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100110; B = 7'b1001000; // Expected: {'P': 7344}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100110; B = 7'b1001000; | Outputs: P=%b | Expected: P=%d",
                 1160,
                 
                 P
                 , 
                 
                 7344
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000010; B = 7'b0110001; // Expected: {'P': 98}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000010; B = 7'b0110001; | Outputs: P=%b | Expected: P=%d",
                 1161,
                 
                 P
                 , 
                 
                 98
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001001; B = 7'b1111011; // Expected: {'P': 8979}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001001; B = 7'b1111011; | Outputs: P=%b | Expected: P=%d",
                 1162,
                 
                 P
                 , 
                 
                 8979
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110101; B = 7'b1111001; // Expected: {'P': 14157}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110101; B = 7'b1111001; | Outputs: P=%b | Expected: P=%d",
                 1163,
                 
                 P
                 , 
                 
                 14157
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000011; B = 7'b0101111; // Expected: {'P': 3149}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000011; B = 7'b0101111; | Outputs: P=%b | Expected: P=%d",
                 1164,
                 
                 P
                 , 
                 
                 3149
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101011; B = 7'b0111111; // Expected: {'P': 6741}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101011; B = 7'b0111111; | Outputs: P=%b | Expected: P=%d",
                 1165,
                 
                 P
                 , 
                 
                 6741
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000000; B = 7'b0111100; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000000; B = 7'b0111100; | Outputs: P=%b | Expected: P=%d",
                 1166,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001111; B = 7'b0010010; // Expected: {'P': 270}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001111; B = 7'b0010010; | Outputs: P=%b | Expected: P=%d",
                 1167,
                 
                 P
                 , 
                 
                 270
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011001; B = 7'b1101000; // Expected: {'P': 9256}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011001; B = 7'b1101000; | Outputs: P=%b | Expected: P=%d",
                 1168,
                 
                 P
                 , 
                 
                 9256
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101000; B = 7'b1101101; // Expected: {'P': 11336}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101000; B = 7'b1101101; | Outputs: P=%b | Expected: P=%d",
                 1169,
                 
                 P
                 , 
                 
                 11336
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100100; B = 7'b1000001; // Expected: {'P': 2340}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100100; B = 7'b1000001; | Outputs: P=%b | Expected: P=%d",
                 1170,
                 
                 P
                 , 
                 
                 2340
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100101; B = 7'b1010100; // Expected: {'P': 8484}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100101; B = 7'b1010100; | Outputs: P=%b | Expected: P=%d",
                 1171,
                 
                 P
                 , 
                 
                 8484
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010000; B = 7'b1000010; // Expected: {'P': 5280}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010000; B = 7'b1000010; | Outputs: P=%b | Expected: P=%d",
                 1172,
                 
                 P
                 , 
                 
                 5280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001100; B = 7'b1010110; // Expected: {'P': 1032}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001100; B = 7'b1010110; | Outputs: P=%b | Expected: P=%d",
                 1173,
                 
                 P
                 , 
                 
                 1032
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000101; B = 7'b0010001; // Expected: {'P': 85}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000101; B = 7'b0010001; | Outputs: P=%b | Expected: P=%d",
                 1174,
                 
                 P
                 , 
                 
                 85
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011011; B = 7'b1000010; // Expected: {'P': 6006}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011011; B = 7'b1000010; | Outputs: P=%b | Expected: P=%d",
                 1175,
                 
                 P
                 , 
                 
                 6006
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010011; B = 7'b1011111; // Expected: {'P': 1805}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010011; B = 7'b1011111; | Outputs: P=%b | Expected: P=%d",
                 1176,
                 
                 P
                 , 
                 
                 1805
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110101; B = 7'b0111110; // Expected: {'P': 7254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110101; B = 7'b0111110; | Outputs: P=%b | Expected: P=%d",
                 1177,
                 
                 P
                 , 
                 
                 7254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111000; B = 7'b1111101; // Expected: {'P': 15000}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111000; B = 7'b1111101; | Outputs: P=%b | Expected: P=%d",
                 1178,
                 
                 P
                 , 
                 
                 15000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101010; B = 7'b1000001; // Expected: {'P': 2730}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101010; B = 7'b1000001; | Outputs: P=%b | Expected: P=%d",
                 1179,
                 
                 P
                 , 
                 
                 2730
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110101; B = 7'b0100000; // Expected: {'P': 3744}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110101; B = 7'b0100000; | Outputs: P=%b | Expected: P=%d",
                 1180,
                 
                 P
                 , 
                 
                 3744
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101100; B = 7'b0101000; // Expected: {'P': 1760}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101100; B = 7'b0101000; | Outputs: P=%b | Expected: P=%d",
                 1181,
                 
                 P
                 , 
                 
                 1760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011000; B = 7'b1010101; // Expected: {'P': 2040}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011000; B = 7'b1010101; | Outputs: P=%b | Expected: P=%d",
                 1182,
                 
                 P
                 , 
                 
                 2040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101011; B = 7'b0011101; // Expected: {'P': 3103}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101011; B = 7'b0011101; | Outputs: P=%b | Expected: P=%d",
                 1183,
                 
                 P
                 , 
                 
                 3103
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110100; B = 7'b0010101; // Expected: {'P': 1092}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110100; B = 7'b0010101; | Outputs: P=%b | Expected: P=%d",
                 1184,
                 
                 P
                 , 
                 
                 1092
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000010; B = 7'b1110101; // Expected: {'P': 7722}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000010; B = 7'b1110101; | Outputs: P=%b | Expected: P=%d",
                 1185,
                 
                 P
                 , 
                 
                 7722
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001110; B = 7'b0101110; // Expected: {'P': 644}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001110; B = 7'b0101110; | Outputs: P=%b | Expected: P=%d",
                 1186,
                 
                 P
                 , 
                 
                 644
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100110; B = 7'b0110111; // Expected: {'P': 2090}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100110; B = 7'b0110111; | Outputs: P=%b | Expected: P=%d",
                 1187,
                 
                 P
                 , 
                 
                 2090
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101001; B = 7'b1110011; // Expected: {'P': 4715}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101001; B = 7'b1110011; | Outputs: P=%b | Expected: P=%d",
                 1188,
                 
                 P
                 , 
                 
                 4715
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110110; B = 7'b1101111; // Expected: {'P': 13098}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110110; B = 7'b1101111; | Outputs: P=%b | Expected: P=%d",
                 1189,
                 
                 P
                 , 
                 
                 13098
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011001; B = 7'b0100111; // Expected: {'P': 3471}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011001; B = 7'b0100111; | Outputs: P=%b | Expected: P=%d",
                 1190,
                 
                 P
                 , 
                 
                 3471
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010010; B = 7'b0110011; // Expected: {'P': 4182}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010010; B = 7'b0110011; | Outputs: P=%b | Expected: P=%d",
                 1191,
                 
                 P
                 , 
                 
                 4182
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111101; B = 7'b0100011; // Expected: {'P': 2135}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111101; B = 7'b0100011; | Outputs: P=%b | Expected: P=%d",
                 1192,
                 
                 P
                 , 
                 
                 2135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110100; B = 7'b0101010; // Expected: {'P': 4872}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110100; B = 7'b0101010; | Outputs: P=%b | Expected: P=%d",
                 1193,
                 
                 P
                 , 
                 
                 4872
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000000; B = 7'b1010000; // Expected: {'P': 5120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000000; B = 7'b1010000; | Outputs: P=%b | Expected: P=%d",
                 1194,
                 
                 P
                 , 
                 
                 5120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111010; B = 7'b0110000; // Expected: {'P': 5856}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111010; B = 7'b0110000; | Outputs: P=%b | Expected: P=%d",
                 1195,
                 
                 P
                 , 
                 
                 5856
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011000; B = 7'b1110001; // Expected: {'P': 9944}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011000; B = 7'b1110001; | Outputs: P=%b | Expected: P=%d",
                 1196,
                 
                 P
                 , 
                 
                 9944
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000011; B = 7'b1001110; // Expected: {'P': 5226}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000011; B = 7'b1001110; | Outputs: P=%b | Expected: P=%d",
                 1197,
                 
                 P
                 , 
                 
                 5226
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101001; B = 7'b0110110; // Expected: {'P': 2214}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101001; B = 7'b0110110; | Outputs: P=%b | Expected: P=%d",
                 1198,
                 
                 P
                 , 
                 
                 2214
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110001; B = 7'b1110110; // Expected: {'P': 13334}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110001; B = 7'b1110110; | Outputs: P=%b | Expected: P=%d",
                 1199,
                 
                 P
                 , 
                 
                 13334
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101010; B = 7'b0110101; // Expected: {'P': 2226}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101010; B = 7'b0110101; | Outputs: P=%b | Expected: P=%d",
                 1200,
                 
                 P
                 , 
                 
                 2226
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100111; B = 7'b0110100; // Expected: {'P': 5356}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100111; B = 7'b0110100; | Outputs: P=%b | Expected: P=%d",
                 1201,
                 
                 P
                 , 
                 
                 5356
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111000; B = 7'b1110100; // Expected: {'P': 6496}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111000; B = 7'b1110100; | Outputs: P=%b | Expected: P=%d",
                 1202,
                 
                 P
                 , 
                 
                 6496
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100101; B = 7'b0101010; // Expected: {'P': 1554}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100101; B = 7'b0101010; | Outputs: P=%b | Expected: P=%d",
                 1203,
                 
                 P
                 , 
                 
                 1554
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001111; B = 7'b1111111; // Expected: {'P': 10033}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001111; B = 7'b1111111; | Outputs: P=%b | Expected: P=%d",
                 1204,
                 
                 P
                 , 
                 
                 10033
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111111; B = 7'b1011111; // Expected: {'P': 5985}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111111; B = 7'b1011111; | Outputs: P=%b | Expected: P=%d",
                 1205,
                 
                 P
                 , 
                 
                 5985
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111010; B = 7'b0101110; // Expected: {'P': 5612}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111010; B = 7'b0101110; | Outputs: P=%b | Expected: P=%d",
                 1206,
                 
                 P
                 , 
                 
                 5612
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010001; B = 7'b0010000; // Expected: {'P': 1296}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010001; B = 7'b0010000; | Outputs: P=%b | Expected: P=%d",
                 1207,
                 
                 P
                 , 
                 
                 1296
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011110; B = 7'b1001101; // Expected: {'P': 2310}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011110; B = 7'b1001101; | Outputs: P=%b | Expected: P=%d",
                 1208,
                 
                 P
                 , 
                 
                 2310
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100001; B = 7'b0010001; // Expected: {'P': 561}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100001; B = 7'b0010001; | Outputs: P=%b | Expected: P=%d",
                 1209,
                 
                 P
                 , 
                 
                 561
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100100; B = 7'b1001100; // Expected: {'P': 7600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100100; B = 7'b1001100; | Outputs: P=%b | Expected: P=%d",
                 1210,
                 
                 P
                 , 
                 
                 7600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010101; B = 7'b1010110; // Expected: {'P': 7310}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010101; B = 7'b1010110; | Outputs: P=%b | Expected: P=%d",
                 1211,
                 
                 P
                 , 
                 
                 7310
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111101; B = 7'b0111100; // Expected: {'P': 3660}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111101; B = 7'b0111100; | Outputs: P=%b | Expected: P=%d",
                 1212,
                 
                 P
                 , 
                 
                 3660
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101101; B = 7'b1011011; // Expected: {'P': 4095}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101101; B = 7'b1011011; | Outputs: P=%b | Expected: P=%d",
                 1213,
                 
                 P
                 , 
                 
                 4095
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010000; B = 7'b1111001; // Expected: {'P': 9680}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010000; B = 7'b1111001; | Outputs: P=%b | Expected: P=%d",
                 1214,
                 
                 P
                 , 
                 
                 9680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100111; B = 7'b0010001; // Expected: {'P': 1751}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100111; B = 7'b0010001; | Outputs: P=%b | Expected: P=%d",
                 1215,
                 
                 P
                 , 
                 
                 1751
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110001; B = 7'b0111100; // Expected: {'P': 6780}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110001; B = 7'b0111100; | Outputs: P=%b | Expected: P=%d",
                 1216,
                 
                 P
                 , 
                 
                 6780
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111101; B = 7'b1100110; // Expected: {'P': 12750}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111101; B = 7'b1100110; | Outputs: P=%b | Expected: P=%d",
                 1217,
                 
                 P
                 , 
                 
                 12750
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011011; B = 7'b0001011; // Expected: {'P': 297}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011011; B = 7'b0001011; | Outputs: P=%b | Expected: P=%d",
                 1218,
                 
                 P
                 , 
                 
                 297
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011110; B = 7'b0111011; // Expected: {'P': 5546}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011110; B = 7'b0111011; | Outputs: P=%b | Expected: P=%d",
                 1219,
                 
                 P
                 , 
                 
                 5546
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010111; B = 7'b0101110; // Expected: {'P': 4002}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010111; B = 7'b0101110; | Outputs: P=%b | Expected: P=%d",
                 1220,
                 
                 P
                 , 
                 
                 4002
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010110; B = 7'b1101000; // Expected: {'P': 8944}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010110; B = 7'b1101000; | Outputs: P=%b | Expected: P=%d",
                 1221,
                 
                 P
                 , 
                 
                 8944
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110001; B = 7'b0010011; // Expected: {'P': 2147}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110001; B = 7'b0010011; | Outputs: P=%b | Expected: P=%d",
                 1222,
                 
                 P
                 , 
                 
                 2147
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011011; B = 7'b0110110; // Expected: {'P': 1458}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011011; B = 7'b0110110; | Outputs: P=%b | Expected: P=%d",
                 1223,
                 
                 P
                 , 
                 
                 1458
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110010; B = 7'b0110010; // Expected: {'P': 5700}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110010; B = 7'b0110010; | Outputs: P=%b | Expected: P=%d",
                 1224,
                 
                 P
                 , 
                 
                 5700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010011; B = 7'b1001010; // Expected: {'P': 1406}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010011; B = 7'b1001010; | Outputs: P=%b | Expected: P=%d",
                 1225,
                 
                 P
                 , 
                 
                 1406
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001111; B = 7'b0111100; // Expected: {'P': 4740}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001111; B = 7'b0111100; | Outputs: P=%b | Expected: P=%d",
                 1226,
                 
                 P
                 , 
                 
                 4740
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011110; B = 7'b0110101; // Expected: {'P': 1590}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011110; B = 7'b0110101; | Outputs: P=%b | Expected: P=%d",
                 1227,
                 
                 P
                 , 
                 
                 1590
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000111; B = 7'b1010101; // Expected: {'P': 6035}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000111; B = 7'b1010101; | Outputs: P=%b | Expected: P=%d",
                 1228,
                 
                 P
                 , 
                 
                 6035
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010110; B = 7'b0001100; // Expected: {'P': 264}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010110; B = 7'b0001100; | Outputs: P=%b | Expected: P=%d",
                 1229,
                 
                 P
                 , 
                 
                 264
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000101; B = 7'b0011000; // Expected: {'P': 120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000101; B = 7'b0011000; | Outputs: P=%b | Expected: P=%d",
                 1230,
                 
                 P
                 , 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111111; B = 7'b0000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111111; B = 7'b0000000; | Outputs: P=%b | Expected: P=%d",
                 1231,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011000; B = 7'b1111111; // Expected: {'P': 11176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011000; B = 7'b1111111; | Outputs: P=%b | Expected: P=%d",
                 1232,
                 
                 P
                 , 
                 
                 11176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000100; B = 7'b1001000; // Expected: {'P': 4896}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000100; B = 7'b1001000; | Outputs: P=%b | Expected: P=%d",
                 1233,
                 
                 P
                 , 
                 
                 4896
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110000; B = 7'b1101000; // Expected: {'P': 4992}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110000; B = 7'b1101000; | Outputs: P=%b | Expected: P=%d",
                 1234,
                 
                 P
                 , 
                 
                 4992
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001100; B = 7'b0011111; // Expected: {'P': 372}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001100; B = 7'b0011111; | Outputs: P=%b | Expected: P=%d",
                 1235,
                 
                 P
                 , 
                 
                 372
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000011; B = 7'b1100100; // Expected: {'P': 6700}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000011; B = 7'b1100100; | Outputs: P=%b | Expected: P=%d",
                 1236,
                 
                 P
                 , 
                 
                 6700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101011; B = 7'b1111000; // Expected: {'P': 5160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101011; B = 7'b1111000; | Outputs: P=%b | Expected: P=%d",
                 1237,
                 
                 P
                 , 
                 
                 5160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111100; B = 7'b0111100; // Expected: {'P': 3600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111100; B = 7'b0111100; | Outputs: P=%b | Expected: P=%d",
                 1238,
                 
                 P
                 , 
                 
                 3600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100001; B = 7'b1101100; // Expected: {'P': 10476}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100001; B = 7'b1101100; | Outputs: P=%b | Expected: P=%d",
                 1239,
                 
                 P
                 , 
                 
                 10476
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010101; B = 7'b1110010; // Expected: {'P': 9690}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010101; B = 7'b1110010; | Outputs: P=%b | Expected: P=%d",
                 1240,
                 
                 P
                 , 
                 
                 9690
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111000; B = 7'b0010010; // Expected: {'P': 1008}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111000; B = 7'b0010010; | Outputs: P=%b | Expected: P=%d",
                 1241,
                 
                 P
                 , 
                 
                 1008
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011000; B = 7'b0010000; // Expected: {'P': 384}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011000; B = 7'b0010000; | Outputs: P=%b | Expected: P=%d",
                 1242,
                 
                 P
                 , 
                 
                 384
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101011; B = 7'b0101101; // Expected: {'P': 4815}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101011; B = 7'b0101101; | Outputs: P=%b | Expected: P=%d",
                 1243,
                 
                 P
                 , 
                 
                 4815
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100101; B = 7'b0001011; // Expected: {'P': 407}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100101; B = 7'b0001011; | Outputs: P=%b | Expected: P=%d",
                 1244,
                 
                 P
                 , 
                 
                 407
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010100; B = 7'b0110001; // Expected: {'P': 980}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010100; B = 7'b0110001; | Outputs: P=%b | Expected: P=%d",
                 1245,
                 
                 P
                 , 
                 
                 980
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100010; B = 7'b0100000; // Expected: {'P': 1088}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100010; B = 7'b0100000; | Outputs: P=%b | Expected: P=%d",
                 1246,
                 
                 P
                 , 
                 
                 1088
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010110; B = 7'b1011010; // Expected: {'P': 1980}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010110; B = 7'b1011010; | Outputs: P=%b | Expected: P=%d",
                 1247,
                 
                 P
                 , 
                 
                 1980
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100001; B = 7'b0000010; // Expected: {'P': 66}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100001; B = 7'b0000010; | Outputs: P=%b | Expected: P=%d",
                 1248,
                 
                 P
                 , 
                 
                 66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111110; B = 7'b1011011; // Expected: {'P': 5642}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111110; B = 7'b1011011; | Outputs: P=%b | Expected: P=%d",
                 1249,
                 
                 P
                 , 
                 
                 5642
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010010; B = 7'b1100100; // Expected: {'P': 1800}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010010; B = 7'b1100100; | Outputs: P=%b | Expected: P=%d",
                 1250,
                 
                 P
                 , 
                 
                 1800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111101; B = 7'b1111000; // Expected: {'P': 15000}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111101; B = 7'b1111000; | Outputs: P=%b | Expected: P=%d",
                 1251,
                 
                 P
                 , 
                 
                 15000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101111; B = 7'b0111100; // Expected: {'P': 6660}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101111; B = 7'b0111100; | Outputs: P=%b | Expected: P=%d",
                 1252,
                 
                 P
                 , 
                 
                 6660
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100000; B = 7'b0110001; // Expected: {'P': 4704}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100000; B = 7'b0110001; | Outputs: P=%b | Expected: P=%d",
                 1253,
                 
                 P
                 , 
                 
                 4704
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111100; B = 7'b0111010; // Expected: {'P': 7192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111100; B = 7'b0111010; | Outputs: P=%b | Expected: P=%d",
                 1254,
                 
                 P
                 , 
                 
                 7192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101011; B = 7'b1100001; // Expected: {'P': 10379}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101011; B = 7'b1100001; | Outputs: P=%b | Expected: P=%d",
                 1255,
                 
                 P
                 , 
                 
                 10379
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111010; B = 7'b0110010; // Expected: {'P': 6100}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111010; B = 7'b0110010; | Outputs: P=%b | Expected: P=%d",
                 1256,
                 
                 P
                 , 
                 
                 6100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111000; B = 7'b1001011; // Expected: {'P': 9000}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111000; B = 7'b1001011; | Outputs: P=%b | Expected: P=%d",
                 1257,
                 
                 P
                 , 
                 
                 9000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000101; B = 7'b0011000; // Expected: {'P': 1656}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000101; B = 7'b0011000; | Outputs: P=%b | Expected: P=%d",
                 1258,
                 
                 P
                 , 
                 
                 1656
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110010; B = 7'b0010100; // Expected: {'P': 1000}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110010; B = 7'b0010100; | Outputs: P=%b | Expected: P=%d",
                 1259,
                 
                 P
                 , 
                 
                 1000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001100; B = 7'b0101111; // Expected: {'P': 564}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001100; B = 7'b0101111; | Outputs: P=%b | Expected: P=%d",
                 1260,
                 
                 P
                 , 
                 
                 564
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101000; B = 7'b0011011; // Expected: {'P': 2808}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101000; B = 7'b0011011; | Outputs: P=%b | Expected: P=%d",
                 1261,
                 
                 P
                 , 
                 
                 2808
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000000; B = 7'b1111110; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000000; B = 7'b1111110; | Outputs: P=%b | Expected: P=%d",
                 1262,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000111; B = 7'b0001111; // Expected: {'P': 105}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000111; B = 7'b0001111; | Outputs: P=%b | Expected: P=%d",
                 1263,
                 
                 P
                 , 
                 
                 105
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000110; B = 7'b1010100; // Expected: {'P': 5880}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000110; B = 7'b1010100; | Outputs: P=%b | Expected: P=%d",
                 1264,
                 
                 P
                 , 
                 
                 5880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011100; B = 7'b1110111; // Expected: {'P': 10948}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011100; B = 7'b1110111; | Outputs: P=%b | Expected: P=%d",
                 1265,
                 
                 P
                 , 
                 
                 10948
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101001; B = 7'b0000011; // Expected: {'P': 123}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101001; B = 7'b0000011; | Outputs: P=%b | Expected: P=%d",
                 1266,
                 
                 P
                 , 
                 
                 123
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011110; B = 7'b0011101; // Expected: {'P': 2726}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011110; B = 7'b0011101; | Outputs: P=%b | Expected: P=%d",
                 1267,
                 
                 P
                 , 
                 
                 2726
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000100; B = 7'b0101101; // Expected: {'P': 180}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000100; B = 7'b0101101; | Outputs: P=%b | Expected: P=%d",
                 1268,
                 
                 P
                 , 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001110; B = 7'b1100111; // Expected: {'P': 8034}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001110; B = 7'b1100111; | Outputs: P=%b | Expected: P=%d",
                 1269,
                 
                 P
                 , 
                 
                 8034
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011001; B = 7'b0110111; // Expected: {'P': 4895}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011001; B = 7'b0110111; | Outputs: P=%b | Expected: P=%d",
                 1270,
                 
                 P
                 , 
                 
                 4895
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101011; B = 7'b0010010; // Expected: {'P': 1926}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101011; B = 7'b0010010; | Outputs: P=%b | Expected: P=%d",
                 1271,
                 
                 P
                 , 
                 
                 1926
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100110; B = 7'b1010010; // Expected: {'P': 3116}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100110; B = 7'b1010010; | Outputs: P=%b | Expected: P=%d",
                 1272,
                 
                 P
                 , 
                 
                 3116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111110; B = 7'b1000011; // Expected: {'P': 8442}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111110; B = 7'b1000011; | Outputs: P=%b | Expected: P=%d",
                 1273,
                 
                 P
                 , 
                 
                 8442
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110001; B = 7'b0111011; // Expected: {'P': 2891}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110001; B = 7'b0111011; | Outputs: P=%b | Expected: P=%d",
                 1274,
                 
                 P
                 , 
                 
                 2891
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010101; B = 7'b1111011; // Expected: {'P': 2583}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010101; B = 7'b1111011; | Outputs: P=%b | Expected: P=%d",
                 1275,
                 
                 P
                 , 
                 
                 2583
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000101; B = 7'b1011000; // Expected: {'P': 6072}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000101; B = 7'b1011000; | Outputs: P=%b | Expected: P=%d",
                 1276,
                 
                 P
                 , 
                 
                 6072
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111110; B = 7'b1011010; // Expected: {'P': 5580}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111110; B = 7'b1011010; | Outputs: P=%b | Expected: P=%d",
                 1277,
                 
                 P
                 , 
                 
                 5580
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010101; B = 7'b0100111; // Expected: {'P': 819}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010101; B = 7'b0100111; | Outputs: P=%b | Expected: P=%d",
                 1278,
                 
                 P
                 , 
                 
                 819
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000110; B = 7'b1100011; // Expected: {'P': 6930}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000110; B = 7'b1100011; | Outputs: P=%b | Expected: P=%d",
                 1279,
                 
                 P
                 , 
                 
                 6930
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010110; B = 7'b0001111; // Expected: {'P': 1290}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010110; B = 7'b0001111; | Outputs: P=%b | Expected: P=%d",
                 1280,
                 
                 P
                 , 
                 
                 1290
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101100; B = 7'b0111010; // Expected: {'P': 6264}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101100; B = 7'b0111010; | Outputs: P=%b | Expected: P=%d",
                 1281,
                 
                 P
                 , 
                 
                 6264
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101100; B = 7'b0110110; // Expected: {'P': 2376}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101100; B = 7'b0110110; | Outputs: P=%b | Expected: P=%d",
                 1282,
                 
                 P
                 , 
                 
                 2376
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001101; B = 7'b0000010; // Expected: {'P': 154}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001101; B = 7'b0000010; | Outputs: P=%b | Expected: P=%d",
                 1283,
                 
                 P
                 , 
                 
                 154
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001001; B = 7'b0110111; // Expected: {'P': 4015}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001001; B = 7'b0110111; | Outputs: P=%b | Expected: P=%d",
                 1284,
                 
                 P
                 , 
                 
                 4015
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101111; B = 7'b1101001; // Expected: {'P': 4935}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101111; B = 7'b1101001; | Outputs: P=%b | Expected: P=%d",
                 1285,
                 
                 P
                 , 
                 
                 4935
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010111; B = 7'b1011000; // Expected: {'P': 2024}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010111; B = 7'b1011000; | Outputs: P=%b | Expected: P=%d",
                 1286,
                 
                 P
                 , 
                 
                 2024
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111011; B = 7'b1110001; // Expected: {'P': 13899}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111011; B = 7'b1110001; | Outputs: P=%b | Expected: P=%d",
                 1287,
                 
                 P
                 , 
                 
                 13899
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100000; B = 7'b1100100; // Expected: {'P': 9600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100000; B = 7'b1100100; | Outputs: P=%b | Expected: P=%d",
                 1288,
                 
                 P
                 , 
                 
                 9600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100100; B = 7'b1000101; // Expected: {'P': 2484}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100100; B = 7'b1000101; | Outputs: P=%b | Expected: P=%d",
                 1289,
                 
                 P
                 , 
                 
                 2484
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011101; B = 7'b0111001; // Expected: {'P': 5301}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011101; B = 7'b0111001; | Outputs: P=%b | Expected: P=%d",
                 1290,
                 
                 P
                 , 
                 
                 5301
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010111; B = 7'b0000010; // Expected: {'P': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010111; B = 7'b0000010; | Outputs: P=%b | Expected: P=%d",
                 1291,
                 
                 P
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001110; B = 7'b1000101; // Expected: {'P': 5382}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001110; B = 7'b1000101; | Outputs: P=%b | Expected: P=%d",
                 1292,
                 
                 P
                 , 
                 
                 5382
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000101; B = 7'b1010110; // Expected: {'P': 5934}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000101; B = 7'b1010110; | Outputs: P=%b | Expected: P=%d",
                 1293,
                 
                 P
                 , 
                 
                 5934
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001111; B = 7'b1100011; // Expected: {'P': 7821}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001111; B = 7'b1100011; | Outputs: P=%b | Expected: P=%d",
                 1294,
                 
                 P
                 , 
                 
                 7821
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101110; B = 7'b1111011; // Expected: {'P': 13530}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101110; B = 7'b1111011; | Outputs: P=%b | Expected: P=%d",
                 1295,
                 
                 P
                 , 
                 
                 13530
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011100; B = 7'b1111100; // Expected: {'P': 11408}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011100; B = 7'b1111100; | Outputs: P=%b | Expected: P=%d",
                 1296,
                 
                 P
                 , 
                 
                 11408
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110011; B = 7'b0101000; // Expected: {'P': 2040}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110011; B = 7'b0101000; | Outputs: P=%b | Expected: P=%d",
                 1297,
                 
                 P
                 , 
                 
                 2040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001001; B = 7'b1011011; // Expected: {'P': 6643}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001001; B = 7'b1011011; | Outputs: P=%b | Expected: P=%d",
                 1298,
                 
                 P
                 , 
                 
                 6643
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001100; B = 7'b1101010; // Expected: {'P': 8056}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001100; B = 7'b1101010; | Outputs: P=%b | Expected: P=%d",
                 1299,
                 
                 P
                 , 
                 
                 8056
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101111; B = 7'b0010000; // Expected: {'P': 752}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101111; B = 7'b0010000; | Outputs: P=%b | Expected: P=%d",
                 1300,
                 
                 P
                 , 
                 
                 752
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100011; B = 7'b1110001; // Expected: {'P': 3955}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100011; B = 7'b1110001; | Outputs: P=%b | Expected: P=%d",
                 1301,
                 
                 P
                 , 
                 
                 3955
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000001; B = 7'b0100101; // Expected: {'P': 2405}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000001; B = 7'b0100101; | Outputs: P=%b | Expected: P=%d",
                 1302,
                 
                 P
                 , 
                 
                 2405
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111000; B = 7'b0010011; // Expected: {'P': 2280}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111000; B = 7'b0010011; | Outputs: P=%b | Expected: P=%d",
                 1303,
                 
                 P
                 , 
                 
                 2280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011111; B = 7'b0101111; // Expected: {'P': 4465}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011111; B = 7'b0101111; | Outputs: P=%b | Expected: P=%d",
                 1304,
                 
                 P
                 , 
                 
                 4465
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111011; B = 7'b1010110; // Expected: {'P': 10578}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111011; B = 7'b1010110; | Outputs: P=%b | Expected: P=%d",
                 1305,
                 
                 P
                 , 
                 
                 10578
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101010; B = 7'b0110101; // Expected: {'P': 5618}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101010; B = 7'b0110101; | Outputs: P=%b | Expected: P=%d",
                 1306,
                 
                 P
                 , 
                 
                 5618
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110010; B = 7'b1101101; // Expected: {'P': 5450}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110010; B = 7'b1101101; | Outputs: P=%b | Expected: P=%d",
                 1307,
                 
                 P
                 , 
                 
                 5450
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010000; B = 7'b1110100; // Expected: {'P': 1856}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010000; B = 7'b1110100; | Outputs: P=%b | Expected: P=%d",
                 1308,
                 
                 P
                 , 
                 
                 1856
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110001; B = 7'b0101001; // Expected: {'P': 4633}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110001; B = 7'b0101001; | Outputs: P=%b | Expected: P=%d",
                 1309,
                 
                 P
                 , 
                 
                 4633
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000111; B = 7'b0100110; // Expected: {'P': 2698}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000111; B = 7'b0100110; | Outputs: P=%b | Expected: P=%d",
                 1310,
                 
                 P
                 , 
                 
                 2698
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100100; B = 7'b1011111; // Expected: {'P': 9500}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100100; B = 7'b1011111; | Outputs: P=%b | Expected: P=%d",
                 1311,
                 
                 P
                 , 
                 
                 9500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001101; B = 7'b0000111; // Expected: {'P': 91}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001101; B = 7'b0000111; | Outputs: P=%b | Expected: P=%d",
                 1312,
                 
                 P
                 , 
                 
                 91
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110001; B = 7'b1011110; // Expected: {'P': 10622}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110001; B = 7'b1011110; | Outputs: P=%b | Expected: P=%d",
                 1313,
                 
                 P
                 , 
                 
                 10622
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010101; B = 7'b1000101; // Expected: {'P': 5865}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010101; B = 7'b1000101; | Outputs: P=%b | Expected: P=%d",
                 1314,
                 
                 P
                 , 
                 
                 5865
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011001; B = 7'b0001000; // Expected: {'P': 712}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011001; B = 7'b0001000; | Outputs: P=%b | Expected: P=%d",
                 1315,
                 
                 P
                 , 
                 
                 712
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010110; B = 7'b0101110; // Expected: {'P': 3956}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010110; B = 7'b0101110; | Outputs: P=%b | Expected: P=%d",
                 1316,
                 
                 P
                 , 
                 
                 3956
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001110; B = 7'b0000010; // Expected: {'P': 156}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001110; B = 7'b0000010; | Outputs: P=%b | Expected: P=%d",
                 1317,
                 
                 P
                 , 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100101; B = 7'b0110101; // Expected: {'P': 1961}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100101; B = 7'b0110101; | Outputs: P=%b | Expected: P=%d",
                 1318,
                 
                 P
                 , 
                 
                 1961
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100100; B = 7'b1010100; // Expected: {'P': 3024}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100100; B = 7'b1010100; | Outputs: P=%b | Expected: P=%d",
                 1319,
                 
                 P
                 , 
                 
                 3024
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001111; B = 7'b0111000; // Expected: {'P': 840}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001111; B = 7'b0111000; | Outputs: P=%b | Expected: P=%d",
                 1320,
                 
                 P
                 , 
                 
                 840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101011; B = 7'b0011001; // Expected: {'P': 2675}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101011; B = 7'b0011001; | Outputs: P=%b | Expected: P=%d",
                 1321,
                 
                 P
                 , 
                 
                 2675
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111101; B = 7'b1001001; // Expected: {'P': 4453}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111101; B = 7'b1001001; | Outputs: P=%b | Expected: P=%d",
                 1322,
                 
                 P
                 , 
                 
                 4453
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001101; B = 7'b1001101; // Expected: {'P': 5929}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001101; B = 7'b1001101; | Outputs: P=%b | Expected: P=%d",
                 1323,
                 
                 P
                 , 
                 
                 5929
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010110; B = 7'b0100110; // Expected: {'P': 3268}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010110; B = 7'b0100110; | Outputs: P=%b | Expected: P=%d",
                 1324,
                 
                 P
                 , 
                 
                 3268
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101100; B = 7'b1110110; // Expected: {'P': 5192}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101100; B = 7'b1110110; | Outputs: P=%b | Expected: P=%d",
                 1325,
                 
                 P
                 , 
                 
                 5192
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111110; B = 7'b1100110; // Expected: {'P': 6324}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111110; B = 7'b1100110; | Outputs: P=%b | Expected: P=%d",
                 1326,
                 
                 P
                 , 
                 
                 6324
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001111; B = 7'b1011110; // Expected: {'P': 7426}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001111; B = 7'b1011110; | Outputs: P=%b | Expected: P=%d",
                 1327,
                 
                 P
                 , 
                 
                 7426
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111001; B = 7'b1001110; // Expected: {'P': 9438}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111001; B = 7'b1001110; | Outputs: P=%b | Expected: P=%d",
                 1328,
                 
                 P
                 , 
                 
                 9438
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011001; B = 7'b0100011; // Expected: {'P': 875}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011001; B = 7'b0100011; | Outputs: P=%b | Expected: P=%d",
                 1329,
                 
                 P
                 , 
                 
                 875
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010011; B = 7'b0111000; // Expected: {'P': 1064}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010011; B = 7'b0111000; | Outputs: P=%b | Expected: P=%d",
                 1330,
                 
                 P
                 , 
                 
                 1064
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110000; B = 7'b1101010; // Expected: {'P': 5088}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110000; B = 7'b1101010; | Outputs: P=%b | Expected: P=%d",
                 1331,
                 
                 P
                 , 
                 
                 5088
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111111; B = 7'b0010100; // Expected: {'P': 2540}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111111; B = 7'b0010100; | Outputs: P=%b | Expected: P=%d",
                 1332,
                 
                 P
                 , 
                 
                 2540
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010010; B = 7'b1111101; // Expected: {'P': 10250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010010; B = 7'b1111101; | Outputs: P=%b | Expected: P=%d",
                 1333,
                 
                 P
                 , 
                 
                 10250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000100; B = 7'b0001100; // Expected: {'P': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000100; B = 7'b0001100; | Outputs: P=%b | Expected: P=%d",
                 1334,
                 
                 P
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010001; B = 7'b0001111; // Expected: {'P': 1215}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010001; B = 7'b0001111; | Outputs: P=%b | Expected: P=%d",
                 1335,
                 
                 P
                 , 
                 
                 1215
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010000; B = 7'b0110001; // Expected: {'P': 784}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010000; B = 7'b0110001; | Outputs: P=%b | Expected: P=%d",
                 1336,
                 
                 P
                 , 
                 
                 784
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001001; B = 7'b0100100; // Expected: {'P': 324}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001001; B = 7'b0100100; | Outputs: P=%b | Expected: P=%d",
                 1337,
                 
                 P
                 , 
                 
                 324
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100101; B = 7'b0000001; // Expected: {'P': 101}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100101; B = 7'b0000001; | Outputs: P=%b | Expected: P=%d",
                 1338,
                 
                 P
                 , 
                 
                 101
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011000; B = 7'b0011011; // Expected: {'P': 648}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011000; B = 7'b0011011; | Outputs: P=%b | Expected: P=%d",
                 1339,
                 
                 P
                 , 
                 
                 648
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011010; B = 7'b0011111; // Expected: {'P': 806}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011010; B = 7'b0011111; | Outputs: P=%b | Expected: P=%d",
                 1340,
                 
                 P
                 , 
                 
                 806
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111100; B = 7'b1011000; // Expected: {'P': 10912}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111100; B = 7'b1011000; | Outputs: P=%b | Expected: P=%d",
                 1341,
                 
                 P
                 , 
                 
                 10912
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010001; B = 7'b0010011; // Expected: {'P': 323}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010001; B = 7'b0010011; | Outputs: P=%b | Expected: P=%d",
                 1342,
                 
                 P
                 , 
                 
                 323
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000100; B = 7'b1111011; // Expected: {'P': 8364}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000100; B = 7'b1111011; | Outputs: P=%b | Expected: P=%d",
                 1343,
                 
                 P
                 , 
                 
                 8364
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011010; B = 7'b0111100; // Expected: {'P': 5400}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011010; B = 7'b0111100; | Outputs: P=%b | Expected: P=%d",
                 1344,
                 
                 P
                 , 
                 
                 5400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001100; B = 7'b1001001; // Expected: {'P': 5548}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001100; B = 7'b1001001; | Outputs: P=%b | Expected: P=%d",
                 1345,
                 
                 P
                 , 
                 
                 5548
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011101; B = 7'b0011100; // Expected: {'P': 812}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011101; B = 7'b0011100; | Outputs: P=%b | Expected: P=%d",
                 1346,
                 
                 P
                 , 
                 
                 812
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111010; B = 7'b0100001; // Expected: {'P': 4026}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111010; B = 7'b0100001; | Outputs: P=%b | Expected: P=%d",
                 1347,
                 
                 P
                 , 
                 
                 4026
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110111; B = 7'b0011100; // Expected: {'P': 3332}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110111; B = 7'b0011100; | Outputs: P=%b | Expected: P=%d",
                 1348,
                 
                 P
                 , 
                 
                 3332
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000010; B = 7'b1001110; // Expected: {'P': 156}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000010; B = 7'b1001110; | Outputs: P=%b | Expected: P=%d",
                 1349,
                 
                 P
                 , 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001011; B = 7'b0110011; // Expected: {'P': 561}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001011; B = 7'b0110011; | Outputs: P=%b | Expected: P=%d",
                 1350,
                 
                 P
                 , 
                 
                 561
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001010; B = 7'b0111000; // Expected: {'P': 560}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001010; B = 7'b0111000; | Outputs: P=%b | Expected: P=%d",
                 1351,
                 
                 P
                 , 
                 
                 560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010100; B = 7'b1100111; // Expected: {'P': 2060}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010100; B = 7'b1100111; | Outputs: P=%b | Expected: P=%d",
                 1352,
                 
                 P
                 , 
                 
                 2060
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110110; B = 7'b1110011; // Expected: {'P': 13570}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110110; B = 7'b1110011; | Outputs: P=%b | Expected: P=%d",
                 1353,
                 
                 P
                 , 
                 
                 13570
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100100; B = 7'b1010111; // Expected: {'P': 8700}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100100; B = 7'b1010111; | Outputs: P=%b | Expected: P=%d",
                 1354,
                 
                 P
                 , 
                 
                 8700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000000; B = 7'b0100100; // Expected: {'P': 2304}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000000; B = 7'b0100100; | Outputs: P=%b | Expected: P=%d",
                 1355,
                 
                 P
                 , 
                 
                 2304
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001001; B = 7'b1110111; // Expected: {'P': 1071}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001001; B = 7'b1110111; | Outputs: P=%b | Expected: P=%d",
                 1356,
                 
                 P
                 , 
                 
                 1071
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111100; B = 7'b1101110; // Expected: {'P': 6600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111100; B = 7'b1101110; | Outputs: P=%b | Expected: P=%d",
                 1357,
                 
                 P
                 , 
                 
                 6600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001101; B = 7'b0111110; // Expected: {'P': 806}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001101; B = 7'b0111110; | Outputs: P=%b | Expected: P=%d",
                 1358,
                 
                 P
                 , 
                 
                 806
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111100; B = 7'b1001011; // Expected: {'P': 4500}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111100; B = 7'b1001011; | Outputs: P=%b | Expected: P=%d",
                 1359,
                 
                 P
                 , 
                 
                 4500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110000; B = 7'b1111111; // Expected: {'P': 6096}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110000; B = 7'b1111111; | Outputs: P=%b | Expected: P=%d",
                 1360,
                 
                 P
                 , 
                 
                 6096
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100100; B = 7'b1011011; // Expected: {'P': 9100}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100100; B = 7'b1011011; | Outputs: P=%b | Expected: P=%d",
                 1361,
                 
                 P
                 , 
                 
                 9100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011001; B = 7'b0001001; // Expected: {'P': 225}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011001; B = 7'b0001001; | Outputs: P=%b | Expected: P=%d",
                 1362,
                 
                 P
                 , 
                 
                 225
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010000; B = 7'b0100000; // Expected: {'P': 2560}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010000; B = 7'b0100000; | Outputs: P=%b | Expected: P=%d",
                 1363,
                 
                 P
                 , 
                 
                 2560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001010; B = 7'b0100011; // Expected: {'P': 2590}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001010; B = 7'b0100011; | Outputs: P=%b | Expected: P=%d",
                 1364,
                 
                 P
                 , 
                 
                 2590
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110011; B = 7'b1010111; // Expected: {'P': 4437}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110011; B = 7'b1010111; | Outputs: P=%b | Expected: P=%d",
                 1365,
                 
                 P
                 , 
                 
                 4437
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110101; B = 7'b0011011; // Expected: {'P': 3159}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110101; B = 7'b0011011; | Outputs: P=%b | Expected: P=%d",
                 1366,
                 
                 P
                 , 
                 
                 3159
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110010; B = 7'b0100111; // Expected: {'P': 4446}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110010; B = 7'b0100111; | Outputs: P=%b | Expected: P=%d",
                 1367,
                 
                 P
                 , 
                 
                 4446
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111101; B = 7'b0101100; // Expected: {'P': 2684}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111101; B = 7'b0101100; | Outputs: P=%b | Expected: P=%d",
                 1368,
                 
                 P
                 , 
                 
                 2684
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001100; B = 7'b0010100; // Expected: {'P': 1520}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001100; B = 7'b0010100; | Outputs: P=%b | Expected: P=%d",
                 1369,
                 
                 P
                 , 
                 
                 1520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000011; B = 7'b1010110; // Expected: {'P': 258}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000011; B = 7'b1010110; | Outputs: P=%b | Expected: P=%d",
                 1370,
                 
                 P
                 , 
                 
                 258
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100100; B = 7'b1100110; // Expected: {'P': 3672}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100100; B = 7'b1100110; | Outputs: P=%b | Expected: P=%d",
                 1371,
                 
                 P
                 , 
                 
                 3672
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110000; B = 7'b0101011; // Expected: {'P': 4816}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110000; B = 7'b0101011; | Outputs: P=%b | Expected: P=%d",
                 1372,
                 
                 P
                 , 
                 
                 4816
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110100; B = 7'b1011100; // Expected: {'P': 4784}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110100; B = 7'b1011100; | Outputs: P=%b | Expected: P=%d",
                 1373,
                 
                 P
                 , 
                 
                 4784
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010100; B = 7'b1111101; // Expected: {'P': 2500}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010100; B = 7'b1111101; | Outputs: P=%b | Expected: P=%d",
                 1374,
                 
                 P
                 , 
                 
                 2500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011010; B = 7'b0111011; // Expected: {'P': 1534}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011010; B = 7'b0111011; | Outputs: P=%b | Expected: P=%d",
                 1375,
                 
                 P
                 , 
                 
                 1534
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100100; B = 7'b1110001; // Expected: {'P': 11300}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100100; B = 7'b1110001; | Outputs: P=%b | Expected: P=%d",
                 1376,
                 
                 P
                 , 
                 
                 11300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110001; B = 7'b0101101; // Expected: {'P': 2205}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110001; B = 7'b0101101; | Outputs: P=%b | Expected: P=%d",
                 1377,
                 
                 P
                 , 
                 
                 2205
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100100; B = 7'b0100111; // Expected: {'P': 1404}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100100; B = 7'b0100111; | Outputs: P=%b | Expected: P=%d",
                 1378,
                 
                 P
                 , 
                 
                 1404
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011100; B = 7'b1000001; // Expected: {'P': 1820}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011100; B = 7'b1000001; | Outputs: P=%b | Expected: P=%d",
                 1379,
                 
                 P
                 , 
                 
                 1820
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100011; B = 7'b0011101; // Expected: {'P': 2871}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100011; B = 7'b0011101; | Outputs: P=%b | Expected: P=%d",
                 1380,
                 
                 P
                 , 
                 
                 2871
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101011; B = 7'b1010000; // Expected: {'P': 8560}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101011; B = 7'b1010000; | Outputs: P=%b | Expected: P=%d",
                 1381,
                 
                 P
                 , 
                 
                 8560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101101; B = 7'b0011001; // Expected: {'P': 2725}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101101; B = 7'b0011001; | Outputs: P=%b | Expected: P=%d",
                 1382,
                 
                 P
                 , 
                 
                 2725
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011011; B = 7'b0101101; // Expected: {'P': 1215}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011011; B = 7'b0101101; | Outputs: P=%b | Expected: P=%d",
                 1383,
                 
                 P
                 , 
                 
                 1215
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101101; B = 7'b1111001; // Expected: {'P': 5445}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101101; B = 7'b1111001; | Outputs: P=%b | Expected: P=%d",
                 1384,
                 
                 P
                 , 
                 
                 5445
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001001; B = 7'b0011001; // Expected: {'P': 1825}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001001; B = 7'b0011001; | Outputs: P=%b | Expected: P=%d",
                 1385,
                 
                 P
                 , 
                 
                 1825
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011100; B = 7'b1011101; // Expected: {'P': 2604}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011100; B = 7'b1011101; | Outputs: P=%b | Expected: P=%d",
                 1386,
                 
                 P
                 , 
                 
                 2604
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111111; B = 7'b0000010; // Expected: {'P': 126}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111111; B = 7'b0000010; | Outputs: P=%b | Expected: P=%d",
                 1387,
                 
                 P
                 , 
                 
                 126
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011000; B = 7'b0101010; // Expected: {'P': 1008}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011000; B = 7'b0101010; | Outputs: P=%b | Expected: P=%d",
                 1388,
                 
                 P
                 , 
                 
                 1008
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011001; B = 7'b0101000; // Expected: {'P': 1000}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011001; B = 7'b0101000; | Outputs: P=%b | Expected: P=%d",
                 1389,
                 
                 P
                 , 
                 
                 1000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000011; B = 7'b1101011; // Expected: {'P': 7169}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000011; B = 7'b1101011; | Outputs: P=%b | Expected: P=%d",
                 1390,
                 
                 P
                 , 
                 
                 7169
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000000; B = 7'b0011000; // Expected: {'P': 1536}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000000; B = 7'b0011000; | Outputs: P=%b | Expected: P=%d",
                 1391,
                 
                 P
                 , 
                 
                 1536
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111011; B = 7'b1111110; // Expected: {'P': 15498}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111011; B = 7'b1111110; | Outputs: P=%b | Expected: P=%d",
                 1392,
                 
                 P
                 , 
                 
                 15498
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100011; B = 7'b1011110; // Expected: {'P': 9306}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100011; B = 7'b1011110; | Outputs: P=%b | Expected: P=%d",
                 1393,
                 
                 P
                 , 
                 
                 9306
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001110; B = 7'b1100010; // Expected: {'P': 1372}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001110; B = 7'b1100010; | Outputs: P=%b | Expected: P=%d",
                 1394,
                 
                 P
                 , 
                 
                 1372
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000110; B = 7'b1101000; // Expected: {'P': 624}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000110; B = 7'b1101000; | Outputs: P=%b | Expected: P=%d",
                 1395,
                 
                 P
                 , 
                 
                 624
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110100; B = 7'b1000001; // Expected: {'P': 7540}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110100; B = 7'b1000001; | Outputs: P=%b | Expected: P=%d",
                 1396,
                 
                 P
                 , 
                 
                 7540
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000110; B = 7'b0010010; // Expected: {'P': 108}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000110; B = 7'b0010010; | Outputs: P=%b | Expected: P=%d",
                 1397,
                 
                 P
                 , 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110010; B = 7'b1001100; // Expected: {'P': 3800}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110010; B = 7'b1001100; | Outputs: P=%b | Expected: P=%d",
                 1398,
                 
                 P
                 , 
                 
                 3800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110010; B = 7'b0000101; // Expected: {'P': 250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110010; B = 7'b0000101; | Outputs: P=%b | Expected: P=%d",
                 1399,
                 
                 P
                 , 
                 
                 250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110111; B = 7'b1101010; // Expected: {'P': 5830}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110111; B = 7'b1101010; | Outputs: P=%b | Expected: P=%d",
                 1400,
                 
                 P
                 , 
                 
                 5830
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111110; B = 7'b1000010; // Expected: {'P': 4092}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111110; B = 7'b1000010; | Outputs: P=%b | Expected: P=%d",
                 1401,
                 
                 P
                 , 
                 
                 4092
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001010; B = 7'b0101101; // Expected: {'P': 450}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001010; B = 7'b0101101; | Outputs: P=%b | Expected: P=%d",
                 1402,
                 
                 P
                 , 
                 
                 450
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000010; B = 7'b0010100; // Expected: {'P': 1320}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000010; B = 7'b0010100; | Outputs: P=%b | Expected: P=%d",
                 1403,
                 
                 P
                 , 
                 
                 1320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010000; B = 7'b0001011; // Expected: {'P': 880}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010000; B = 7'b0001011; | Outputs: P=%b | Expected: P=%d",
                 1404,
                 
                 P
                 , 
                 
                 880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110011; B = 7'b0011010; // Expected: {'P': 1326}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110011; B = 7'b0011010; | Outputs: P=%b | Expected: P=%d",
                 1405,
                 
                 P
                 , 
                 
                 1326
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111000; B = 7'b1001100; // Expected: {'P': 4256}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111000; B = 7'b1001100; | Outputs: P=%b | Expected: P=%d",
                 1406,
                 
                 P
                 , 
                 
                 4256
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111000; B = 7'b0001011; // Expected: {'P': 1320}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111000; B = 7'b0001011; | Outputs: P=%b | Expected: P=%d",
                 1407,
                 
                 P
                 , 
                 
                 1320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100000; B = 7'b1101001; // Expected: {'P': 10080}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100000; B = 7'b1101001; | Outputs: P=%b | Expected: P=%d",
                 1408,
                 
                 P
                 , 
                 
                 10080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001001; B = 7'b0011110; // Expected: {'P': 270}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001001; B = 7'b0011110; | Outputs: P=%b | Expected: P=%d",
                 1409,
                 
                 P
                 , 
                 
                 270
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101100; B = 7'b0100100; // Expected: {'P': 3888}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101100; B = 7'b0100100; | Outputs: P=%b | Expected: P=%d",
                 1410,
                 
                 P
                 , 
                 
                 3888
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000110; B = 7'b0110111; // Expected: {'P': 330}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000110; B = 7'b0110111; | Outputs: P=%b | Expected: P=%d",
                 1411,
                 
                 P
                 , 
                 
                 330
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011110; B = 7'b0010101; // Expected: {'P': 1974}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011110; B = 7'b0010101; | Outputs: P=%b | Expected: P=%d",
                 1412,
                 
                 P
                 , 
                 
                 1974
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000001; B = 7'b0010111; // Expected: {'P': 1495}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000001; B = 7'b0010111; | Outputs: P=%b | Expected: P=%d",
                 1413,
                 
                 P
                 , 
                 
                 1495
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110000; B = 7'b0110111; // Expected: {'P': 2640}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110000; B = 7'b0110111; | Outputs: P=%b | Expected: P=%d",
                 1414,
                 
                 P
                 , 
                 
                 2640
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010011; B = 7'b0011111; // Expected: {'P': 589}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010011; B = 7'b0011111; | Outputs: P=%b | Expected: P=%d",
                 1415,
                 
                 P
                 , 
                 
                 589
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100101; B = 7'b0000101; // Expected: {'P': 185}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100101; B = 7'b0000101; | Outputs: P=%b | Expected: P=%d",
                 1416,
                 
                 P
                 , 
                 
                 185
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001101; B = 7'b0110001; // Expected: {'P': 3773}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001101; B = 7'b0110001; | Outputs: P=%b | Expected: P=%d",
                 1417,
                 
                 P
                 , 
                 
                 3773
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110110; B = 7'b0101010; // Expected: {'P': 4956}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110110; B = 7'b0101010; | Outputs: P=%b | Expected: P=%d",
                 1418,
                 
                 P
                 , 
                 
                 4956
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001000; B = 7'b0001001; // Expected: {'P': 72}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001000; B = 7'b0001001; | Outputs: P=%b | Expected: P=%d",
                 1419,
                 
                 P
                 , 
                 
                 72
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011001; B = 7'b1111001; // Expected: {'P': 10769}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011001; B = 7'b1111001; | Outputs: P=%b | Expected: P=%d",
                 1420,
                 
                 P
                 , 
                 
                 10769
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101011; B = 7'b1001110; // Expected: {'P': 8346}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101011; B = 7'b1001110; | Outputs: P=%b | Expected: P=%d",
                 1421,
                 
                 P
                 , 
                 
                 8346
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001011; B = 7'b1101101; // Expected: {'P': 1199}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001011; B = 7'b1101101; | Outputs: P=%b | Expected: P=%d",
                 1422,
                 
                 P
                 , 
                 
                 1199
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001100; B = 7'b1100000; // Expected: {'P': 1152}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001100; B = 7'b1100000; | Outputs: P=%b | Expected: P=%d",
                 1423,
                 
                 P
                 , 
                 
                 1152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011010; B = 7'b1000010; // Expected: {'P': 5940}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011010; B = 7'b1000010; | Outputs: P=%b | Expected: P=%d",
                 1424,
                 
                 P
                 , 
                 
                 5940
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111011; B = 7'b1100101; // Expected: {'P': 5959}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111011; B = 7'b1100101; | Outputs: P=%b | Expected: P=%d",
                 1425,
                 
                 P
                 , 
                 
                 5959
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100011; B = 7'b1110101; // Expected: {'P': 4095}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100011; B = 7'b1110101; | Outputs: P=%b | Expected: P=%d",
                 1426,
                 
                 P
                 , 
                 
                 4095
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101011; B = 7'b0111011; // Expected: {'P': 2537}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101011; B = 7'b0111011; | Outputs: P=%b | Expected: P=%d",
                 1427,
                 
                 P
                 , 
                 
                 2537
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110010; B = 7'b1011010; // Expected: {'P': 4500}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110010; B = 7'b1011010; | Outputs: P=%b | Expected: P=%d",
                 1428,
                 
                 P
                 , 
                 
                 4500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011100; B = 7'b1110110; // Expected: {'P': 10856}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011100; B = 7'b1110110; | Outputs: P=%b | Expected: P=%d",
                 1429,
                 
                 P
                 , 
                 
                 10856
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010010; B = 7'b0101010; // Expected: {'P': 756}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010010; B = 7'b0101010; | Outputs: P=%b | Expected: P=%d",
                 1430,
                 
                 P
                 , 
                 
                 756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110101; B = 7'b1001011; // Expected: {'P': 3975}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110101; B = 7'b1001011; | Outputs: P=%b | Expected: P=%d",
                 1431,
                 
                 P
                 , 
                 
                 3975
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100110; B = 7'b0010111; // Expected: {'P': 2346}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100110; B = 7'b0010111; | Outputs: P=%b | Expected: P=%d",
                 1432,
                 
                 P
                 , 
                 
                 2346
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001111; B = 7'b0011000; // Expected: {'P': 1896}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001111; B = 7'b0011000; | Outputs: P=%b | Expected: P=%d",
                 1433,
                 
                 P
                 , 
                 
                 1896
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011011; B = 7'b0000011; // Expected: {'P': 81}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011011; B = 7'b0000011; | Outputs: P=%b | Expected: P=%d",
                 1434,
                 
                 P
                 , 
                 
                 81
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101011; B = 7'b0010101; // Expected: {'P': 2247}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101011; B = 7'b0010101; | Outputs: P=%b | Expected: P=%d",
                 1435,
                 
                 P
                 , 
                 
                 2247
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111111; B = 7'b0001101; // Expected: {'P': 1651}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111111; B = 7'b0001101; | Outputs: P=%b | Expected: P=%d",
                 1436,
                 
                 P
                 , 
                 
                 1651
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011011; B = 7'b1100000; // Expected: {'P': 2592}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011011; B = 7'b1100000; | Outputs: P=%b | Expected: P=%d",
                 1437,
                 
                 P
                 , 
                 
                 2592
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111010; B = 7'b0011000; // Expected: {'P': 2928}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111010; B = 7'b0011000; | Outputs: P=%b | Expected: P=%d",
                 1438,
                 
                 P
                 , 
                 
                 2928
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100011; B = 7'b1100000; // Expected: {'P': 3360}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100011; B = 7'b1100000; | Outputs: P=%b | Expected: P=%d",
                 1439,
                 
                 P
                 , 
                 
                 3360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100010; B = 7'b1000010; // Expected: {'P': 6468}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100010; B = 7'b1000010; | Outputs: P=%b | Expected: P=%d",
                 1440,
                 
                 P
                 , 
                 
                 6468
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011000; B = 7'b1101101; // Expected: {'P': 2616}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011000; B = 7'b1101101; | Outputs: P=%b | Expected: P=%d",
                 1441,
                 
                 P
                 , 
                 
                 2616
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100001; B = 7'b1011110; // Expected: {'P': 3102}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100001; B = 7'b1011110; | Outputs: P=%b | Expected: P=%d",
                 1442,
                 
                 P
                 , 
                 
                 3102
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101001; B = 7'b1111110; // Expected: {'P': 5166}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101001; B = 7'b1111110; | Outputs: P=%b | Expected: P=%d",
                 1443,
                 
                 P
                 , 
                 
                 5166
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110000; B = 7'b0001110; // Expected: {'P': 1568}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110000; B = 7'b0001110; | Outputs: P=%b | Expected: P=%d",
                 1444,
                 
                 P
                 , 
                 
                 1568
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110000; B = 7'b1011101; // Expected: {'P': 10416}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110000; B = 7'b1011101; | Outputs: P=%b | Expected: P=%d",
                 1445,
                 
                 P
                 , 
                 
                 10416
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101011; B = 7'b1011001; // Expected: {'P': 3827}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101011; B = 7'b1011001; | Outputs: P=%b | Expected: P=%d",
                 1446,
                 
                 P
                 , 
                 
                 3827
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100010; B = 7'b0111110; // Expected: {'P': 6076}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100010; B = 7'b0111110; | Outputs: P=%b | Expected: P=%d",
                 1447,
                 
                 P
                 , 
                 
                 6076
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110000; B = 7'b0100010; // Expected: {'P': 3808}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110000; B = 7'b0100010; | Outputs: P=%b | Expected: P=%d",
                 1448,
                 
                 P
                 , 
                 
                 3808
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000000; B = 7'b0101000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000000; B = 7'b0101000; | Outputs: P=%b | Expected: P=%d",
                 1449,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110000; B = 7'b1000010; // Expected: {'P': 3168}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110000; B = 7'b1000010; | Outputs: P=%b | Expected: P=%d",
                 1450,
                 
                 P
                 , 
                 
                 3168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011101; B = 7'b1100100; // Expected: {'P': 9300}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011101; B = 7'b1100100; | Outputs: P=%b | Expected: P=%d",
                 1451,
                 
                 P
                 , 
                 
                 9300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010110; B = 7'b0100010; // Expected: {'P': 2924}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010110; B = 7'b0100010; | Outputs: P=%b | Expected: P=%d",
                 1452,
                 
                 P
                 , 
                 
                 2924
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111011; B = 7'b0111100; // Expected: {'P': 7380}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111011; B = 7'b0111100; | Outputs: P=%b | Expected: P=%d",
                 1453,
                 
                 P
                 , 
                 
                 7380
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000101; B = 7'b0011010; // Expected: {'P': 1794}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000101; B = 7'b0011010; | Outputs: P=%b | Expected: P=%d",
                 1454,
                 
                 P
                 , 
                 
                 1794
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100001; B = 7'b1111110; // Expected: {'P': 12222}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100001; B = 7'b1111110; | Outputs: P=%b | Expected: P=%d",
                 1455,
                 
                 P
                 , 
                 
                 12222
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100001; B = 7'b1110011; // Expected: {'P': 11155}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100001; B = 7'b1110011; | Outputs: P=%b | Expected: P=%d",
                 1456,
                 
                 P
                 , 
                 
                 11155
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011010; B = 7'b0101100; // Expected: {'P': 3960}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011010; B = 7'b0101100; | Outputs: P=%b | Expected: P=%d",
                 1457,
                 
                 P
                 , 
                 
                 3960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101011; B = 7'b1101010; // Expected: {'P': 11342}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101011; B = 7'b1101010; | Outputs: P=%b | Expected: P=%d",
                 1458,
                 
                 P
                 , 
                 
                 11342
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110011; B = 7'b1110111; // Expected: {'P': 6069}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110011; B = 7'b1110111; | Outputs: P=%b | Expected: P=%d",
                 1459,
                 
                 P
                 , 
                 
                 6069
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011111; B = 7'b0000101; // Expected: {'P': 155}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011111; B = 7'b0000101; | Outputs: P=%b | Expected: P=%d",
                 1460,
                 
                 P
                 , 
                 
                 155
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100010; B = 7'b1111001; // Expected: {'P': 11858}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100010; B = 7'b1111001; | Outputs: P=%b | Expected: P=%d",
                 1461,
                 
                 P
                 , 
                 
                 11858
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010000; B = 7'b1110000; // Expected: {'P': 8960}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010000; B = 7'b1110000; | Outputs: P=%b | Expected: P=%d",
                 1462,
                 
                 P
                 , 
                 
                 8960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100001; B = 7'b1110001; // Expected: {'P': 3729}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100001; B = 7'b1110001; | Outputs: P=%b | Expected: P=%d",
                 1463,
                 
                 P
                 , 
                 
                 3729
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010000; B = 7'b1011001; // Expected: {'P': 7120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010000; B = 7'b1011001; | Outputs: P=%b | Expected: P=%d",
                 1464,
                 
                 P
                 , 
                 
                 7120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001110; B = 7'b1011110; // Expected: {'P': 1316}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001110; B = 7'b1011110; | Outputs: P=%b | Expected: P=%d",
                 1465,
                 
                 P
                 , 
                 
                 1316
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110111; B = 7'b1001011; // Expected: {'P': 8925}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110111; B = 7'b1001011; | Outputs: P=%b | Expected: P=%d",
                 1466,
                 
                 P
                 , 
                 
                 8925
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000110; B = 7'b0011000; // Expected: {'P': 144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000110; B = 7'b0011000; | Outputs: P=%b | Expected: P=%d",
                 1467,
                 
                 P
                 , 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001001; B = 7'b1101100; // Expected: {'P': 7884}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001001; B = 7'b1101100; | Outputs: P=%b | Expected: P=%d",
                 1468,
                 
                 P
                 , 
                 
                 7884
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001000; B = 7'b1010000; // Expected: {'P': 5760}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001000; B = 7'b1010000; | Outputs: P=%b | Expected: P=%d",
                 1469,
                 
                 P
                 , 
                 
                 5760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001001; B = 7'b0010010; // Expected: {'P': 1314}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001001; B = 7'b0010010; | Outputs: P=%b | Expected: P=%d",
                 1470,
                 
                 P
                 , 
                 
                 1314
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100101; B = 7'b1110101; // Expected: {'P': 11817}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100101; B = 7'b1110101; | Outputs: P=%b | Expected: P=%d",
                 1471,
                 
                 P
                 , 
                 
                 11817
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001111; B = 7'b1110100; // Expected: {'P': 1740}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001111; B = 7'b1110100; | Outputs: P=%b | Expected: P=%d",
                 1472,
                 
                 P
                 , 
                 
                 1740
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010100; B = 7'b1010000; // Expected: {'P': 6720}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010100; B = 7'b1010000; | Outputs: P=%b | Expected: P=%d",
                 1473,
                 
                 P
                 , 
                 
                 6720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010111; B = 7'b0101010; // Expected: {'P': 966}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010111; B = 7'b0101010; | Outputs: P=%b | Expected: P=%d",
                 1474,
                 
                 P
                 , 
                 
                 966
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010001; B = 7'b0001011; // Expected: {'P': 891}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010001; B = 7'b0001011; | Outputs: P=%b | Expected: P=%d",
                 1475,
                 
                 P
                 , 
                 
                 891
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110100; B = 7'b0100011; // Expected: {'P': 1820}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110100; B = 7'b0100011; | Outputs: P=%b | Expected: P=%d",
                 1476,
                 
                 P
                 , 
                 
                 1820
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000011; B = 7'b0110000; // Expected: {'P': 144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000011; B = 7'b0110000; | Outputs: P=%b | Expected: P=%d",
                 1477,
                 
                 P
                 , 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110111; B = 7'b0100111; // Expected: {'P': 2145}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110111; B = 7'b0100111; | Outputs: P=%b | Expected: P=%d",
                 1478,
                 
                 P
                 , 
                 
                 2145
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010101; B = 7'b0111000; // Expected: {'P': 1176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010101; B = 7'b0111000; | Outputs: P=%b | Expected: P=%d",
                 1479,
                 
                 P
                 , 
                 
                 1176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001011; B = 7'b1010100; // Expected: {'P': 924}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001011; B = 7'b1010100; | Outputs: P=%b | Expected: P=%d",
                 1480,
                 
                 P
                 , 
                 
                 924
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010100; B = 7'b0001001; // Expected: {'P': 180}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010100; B = 7'b0001001; | Outputs: P=%b | Expected: P=%d",
                 1481,
                 
                 P
                 , 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000011; B = 7'b0010110; // Expected: {'P': 66}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000011; B = 7'b0010110; | Outputs: P=%b | Expected: P=%d",
                 1482,
                 
                 P
                 , 
                 
                 66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111011; B = 7'b0011000; // Expected: {'P': 1416}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111011; B = 7'b0011000; | Outputs: P=%b | Expected: P=%d",
                 1483,
                 
                 P
                 , 
                 
                 1416
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011111; B = 7'b1101000; // Expected: {'P': 3224}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011111; B = 7'b1101000; | Outputs: P=%b | Expected: P=%d",
                 1484,
                 
                 P
                 , 
                 
                 3224
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011101; B = 7'b0100100; // Expected: {'P': 3348}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011101; B = 7'b0100100; | Outputs: P=%b | Expected: P=%d",
                 1485,
                 
                 P
                 , 
                 
                 3348
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100010; B = 7'b1000011; // Expected: {'P': 2278}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100010; B = 7'b1000011; | Outputs: P=%b | Expected: P=%d",
                 1486,
                 
                 P
                 , 
                 
                 2278
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011000; B = 7'b0111111; // Expected: {'P': 5544}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011000; B = 7'b0111111; | Outputs: P=%b | Expected: P=%d",
                 1487,
                 
                 P
                 , 
                 
                 5544
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001010; B = 7'b0000111; // Expected: {'P': 518}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001010; B = 7'b0000111; | Outputs: P=%b | Expected: P=%d",
                 1488,
                 
                 P
                 , 
                 
                 518
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110011; B = 7'b0100110; // Expected: {'P': 1938}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110011; B = 7'b0100110; | Outputs: P=%b | Expected: P=%d",
                 1489,
                 
                 P
                 , 
                 
                 1938
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000001; B = 7'b0111001; // Expected: {'P': 3705}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000001; B = 7'b0111001; | Outputs: P=%b | Expected: P=%d",
                 1490,
                 
                 P
                 , 
                 
                 3705
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000110; B = 7'b1100111; // Expected: {'P': 7210}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000110; B = 7'b1100111; | Outputs: P=%b | Expected: P=%d",
                 1491,
                 
                 P
                 , 
                 
                 7210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001111; B = 7'b1001101; // Expected: {'P': 6083}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001111; B = 7'b1001101; | Outputs: P=%b | Expected: P=%d",
                 1492,
                 
                 P
                 , 
                 
                 6083
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101011; B = 7'b1001101; // Expected: {'P': 3311}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101011; B = 7'b1001101; | Outputs: P=%b | Expected: P=%d",
                 1493,
                 
                 P
                 , 
                 
                 3311
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111011; B = 7'b1010110; // Expected: {'P': 5074}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111011; B = 7'b1010110; | Outputs: P=%b | Expected: P=%d",
                 1494,
                 
                 P
                 , 
                 
                 5074
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100110; B = 7'b1001011; // Expected: {'P': 2850}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100110; B = 7'b1001011; | Outputs: P=%b | Expected: P=%d",
                 1495,
                 
                 P
                 , 
                 
                 2850
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001101; B = 7'b1011001; // Expected: {'P': 1157}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001101; B = 7'b1011001; | Outputs: P=%b | Expected: P=%d",
                 1496,
                 
                 P
                 , 
                 
                 1157
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010100; B = 7'b0110101; // Expected: {'P': 1060}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010100; B = 7'b0110101; | Outputs: P=%b | Expected: P=%d",
                 1497,
                 
                 P
                 , 
                 
                 1060
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001010; B = 7'b0010101; // Expected: {'P': 210}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001010; B = 7'b0010101; | Outputs: P=%b | Expected: P=%d",
                 1498,
                 
                 P
                 , 
                 
                 210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101011; B = 7'b1100010; // Expected: {'P': 10486}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101011; B = 7'b1100010; | Outputs: P=%b | Expected: P=%d",
                 1499,
                 
                 P
                 , 
                 
                 10486
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110100; B = 7'b1100100; // Expected: {'P': 11600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110100; B = 7'b1100100; | Outputs: P=%b | Expected: P=%d",
                 1500,
                 
                 P
                 , 
                 
                 11600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101001; B = 7'b1010111; // Expected: {'P': 9135}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101001; B = 7'b1010111; | Outputs: P=%b | Expected: P=%d",
                 1501,
                 
                 P
                 , 
                 
                 9135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111011; B = 7'b0100110; // Expected: {'P': 2242}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111011; B = 7'b0100110; | Outputs: P=%b | Expected: P=%d",
                 1502,
                 
                 P
                 , 
                 
                 2242
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001000; B = 7'b0101011; // Expected: {'P': 344}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001000; B = 7'b0101011; | Outputs: P=%b | Expected: P=%d",
                 1503,
                 
                 P
                 , 
                 
                 344
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101010; B = 7'b1111110; // Expected: {'P': 13356}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101010; B = 7'b1111110; | Outputs: P=%b | Expected: P=%d",
                 1504,
                 
                 P
                 , 
                 
                 13356
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010111; B = 7'b1010111; // Expected: {'P': 2001}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010111; B = 7'b1010111; | Outputs: P=%b | Expected: P=%d",
                 1505,
                 
                 P
                 , 
                 
                 2001
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010001; B = 7'b1111110; // Expected: {'P': 10206}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010001; B = 7'b1111110; | Outputs: P=%b | Expected: P=%d",
                 1506,
                 
                 P
                 , 
                 
                 10206
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001110; B = 7'b0000001; // Expected: {'P': 78}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001110; B = 7'b0000001; | Outputs: P=%b | Expected: P=%d",
                 1507,
                 
                 P
                 , 
                 
                 78
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100001; B = 7'b1101101; // Expected: {'P': 3597}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100001; B = 7'b1101101; | Outputs: P=%b | Expected: P=%d",
                 1508,
                 
                 P
                 , 
                 
                 3597
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010110; B = 7'b1100000; // Expected: {'P': 8256}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010110; B = 7'b1100000; | Outputs: P=%b | Expected: P=%d",
                 1509,
                 
                 P
                 , 
                 
                 8256
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101011; B = 7'b1000111; // Expected: {'P': 3053}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101011; B = 7'b1000111; | Outputs: P=%b | Expected: P=%d",
                 1510,
                 
                 P
                 , 
                 
                 3053
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110110; B = 7'b0100100; // Expected: {'P': 4248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110110; B = 7'b0100100; | Outputs: P=%b | Expected: P=%d",
                 1511,
                 
                 P
                 , 
                 
                 4248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111110; B = 7'b0010000; // Expected: {'P': 2016}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111110; B = 7'b0010000; | Outputs: P=%b | Expected: P=%d",
                 1512,
                 
                 P
                 , 
                 
                 2016
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110010; B = 7'b0001000; // Expected: {'P': 400}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110010; B = 7'b0001000; | Outputs: P=%b | Expected: P=%d",
                 1513,
                 
                 P
                 , 
                 
                 400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001000; B = 7'b0100001; // Expected: {'P': 2376}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001000; B = 7'b0100001; | Outputs: P=%b | Expected: P=%d",
                 1514,
                 
                 P
                 , 
                 
                 2376
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001101; B = 7'b1011101; // Expected: {'P': 1209}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001101; B = 7'b1011101; | Outputs: P=%b | Expected: P=%d",
                 1515,
                 
                 P
                 , 
                 
                 1209
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101011; B = 7'b1101001; // Expected: {'P': 4515}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101011; B = 7'b1101001; | Outputs: P=%b | Expected: P=%d",
                 1516,
                 
                 P
                 , 
                 
                 4515
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000111; B = 7'b1111101; // Expected: {'P': 8875}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000111; B = 7'b1111101; | Outputs: P=%b | Expected: P=%d",
                 1517,
                 
                 P
                 , 
                 
                 8875
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001001; B = 7'b1101101; // Expected: {'P': 981}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001001; B = 7'b1101101; | Outputs: P=%b | Expected: P=%d",
                 1518,
                 
                 P
                 , 
                 
                 981
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000011; B = 7'b1100110; // Expected: {'P': 6834}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000011; B = 7'b1100110; | Outputs: P=%b | Expected: P=%d",
                 1519,
                 
                 P
                 , 
                 
                 6834
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001001; B = 7'b0001010; // Expected: {'P': 730}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001001; B = 7'b0001010; | Outputs: P=%b | Expected: P=%d",
                 1520,
                 
                 P
                 , 
                 
                 730
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110011; B = 7'b0101111; // Expected: {'P': 2397}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110011; B = 7'b0101111; | Outputs: P=%b | Expected: P=%d",
                 1521,
                 
                 P
                 , 
                 
                 2397
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001111; B = 7'b1100001; // Expected: {'P': 1455}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001111; B = 7'b1100001; | Outputs: P=%b | Expected: P=%d",
                 1522,
                 
                 P
                 , 
                 
                 1455
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001001; B = 7'b0001101; // Expected: {'P': 949}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001001; B = 7'b0001101; | Outputs: P=%b | Expected: P=%d",
                 1523,
                 
                 P
                 , 
                 
                 949
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101100; B = 7'b1101010; // Expected: {'P': 4664}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101100; B = 7'b1101010; | Outputs: P=%b | Expected: P=%d",
                 1524,
                 
                 P
                 , 
                 
                 4664
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010010; B = 7'b0011101; // Expected: {'P': 2378}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010010; B = 7'b0011101; | Outputs: P=%b | Expected: P=%d",
                 1525,
                 
                 P
                 , 
                 
                 2378
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011010; B = 7'b0101110; // Expected: {'P': 1196}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011010; B = 7'b0101110; | Outputs: P=%b | Expected: P=%d",
                 1526,
                 
                 P
                 , 
                 
                 1196
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101110; B = 7'b0100011; // Expected: {'P': 1610}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101110; B = 7'b0100011; | Outputs: P=%b | Expected: P=%d",
                 1527,
                 
                 P
                 , 
                 
                 1610
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100011; B = 7'b0010001; // Expected: {'P': 595}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100011; B = 7'b0010001; | Outputs: P=%b | Expected: P=%d",
                 1528,
                 
                 P
                 , 
                 
                 595
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010111; B = 7'b1100000; // Expected: {'P': 2208}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010111; B = 7'b1100000; | Outputs: P=%b | Expected: P=%d",
                 1529,
                 
                 P
                 , 
                 
                 2208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010100; B = 7'b1100110; // Expected: {'P': 8568}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010100; B = 7'b1100110; | Outputs: P=%b | Expected: P=%d",
                 1530,
                 
                 P
                 , 
                 
                 8568
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000001; B = 7'b0001000; // Expected: {'P': 8}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000001; B = 7'b0001000; | Outputs: P=%b | Expected: P=%d",
                 1531,
                 
                 P
                 , 
                 
                 8
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101000; B = 7'b1111011; // Expected: {'P': 4920}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101000; B = 7'b1111011; | Outputs: P=%b | Expected: P=%d",
                 1532,
                 
                 P
                 , 
                 
                 4920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101110; B = 7'b0010010; // Expected: {'P': 828}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101110; B = 7'b0010010; | Outputs: P=%b | Expected: P=%d",
                 1533,
                 
                 P
                 , 
                 
                 828
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011011; B = 7'b0110000; // Expected: {'P': 1296}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011011; B = 7'b0110000; | Outputs: P=%b | Expected: P=%d",
                 1534,
                 
                 P
                 , 
                 
                 1296
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101101; B = 7'b0010011; // Expected: {'P': 855}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101101; B = 7'b0010011; | Outputs: P=%b | Expected: P=%d",
                 1535,
                 
                 P
                 , 
                 
                 855
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010100; B = 7'b0000010; // Expected: {'P': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010100; B = 7'b0000010; | Outputs: P=%b | Expected: P=%d",
                 1536,
                 
                 P
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000111; B = 7'b0001001; // Expected: {'P': 63}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000111; B = 7'b0001001; | Outputs: P=%b | Expected: P=%d",
                 1537,
                 
                 P
                 , 
                 
                 63
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100100; B = 7'b0101011; // Expected: {'P': 4300}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100100; B = 7'b0101011; | Outputs: P=%b | Expected: P=%d",
                 1538,
                 
                 P
                 , 
                 
                 4300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000000; B = 7'b0100111; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000000; B = 7'b0100111; | Outputs: P=%b | Expected: P=%d",
                 1539,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011100; B = 7'b1111111; // Expected: {'P': 11684}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011100; B = 7'b1111111; | Outputs: P=%b | Expected: P=%d",
                 1540,
                 
                 P
                 , 
                 
                 11684
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001010; B = 7'b0010001; // Expected: {'P': 170}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001010; B = 7'b0010001; | Outputs: P=%b | Expected: P=%d",
                 1541,
                 
                 P
                 , 
                 
                 170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000000; B = 7'b0111000; // Expected: {'P': 3584}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000000; B = 7'b0111000; | Outputs: P=%b | Expected: P=%d",
                 1542,
                 
                 P
                 , 
                 
                 3584
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000111; B = 7'b1100100; // Expected: {'P': 700}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000111; B = 7'b1100100; | Outputs: P=%b | Expected: P=%d",
                 1543,
                 
                 P
                 , 
                 
                 700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011101; B = 7'b1000100; // Expected: {'P': 6324}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011101; B = 7'b1000100; | Outputs: P=%b | Expected: P=%d",
                 1544,
                 
                 P
                 , 
                 
                 6324
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000100; B = 7'b1101110; // Expected: {'P': 440}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000100; B = 7'b1101110; | Outputs: P=%b | Expected: P=%d",
                 1545,
                 
                 P
                 , 
                 
                 440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000011; B = 7'b1101110; // Expected: {'P': 7370}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000011; B = 7'b1101110; | Outputs: P=%b | Expected: P=%d",
                 1546,
                 
                 P
                 , 
                 
                 7370
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000000; B = 7'b1111101; // Expected: {'P': 8000}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000000; B = 7'b1111101; | Outputs: P=%b | Expected: P=%d",
                 1547,
                 
                 P
                 , 
                 
                 8000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010010; B = 7'b1100001; // Expected: {'P': 7954}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010010; B = 7'b1100001; | Outputs: P=%b | Expected: P=%d",
                 1548,
                 
                 P
                 , 
                 
                 7954
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101100; B = 7'b1100001; // Expected: {'P': 4268}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101100; B = 7'b1100001; | Outputs: P=%b | Expected: P=%d",
                 1549,
                 
                 P
                 , 
                 
                 4268
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110110; B = 7'b1111011; // Expected: {'P': 6642}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110110; B = 7'b1111011; | Outputs: P=%b | Expected: P=%d",
                 1550,
                 
                 P
                 , 
                 
                 6642
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001101; B = 7'b1010000; // Expected: {'P': 1040}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001101; B = 7'b1010000; | Outputs: P=%b | Expected: P=%d",
                 1551,
                 
                 P
                 , 
                 
                 1040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001010; B = 7'b1100110; // Expected: {'P': 7548}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001010; B = 7'b1100110; | Outputs: P=%b | Expected: P=%d",
                 1552,
                 
                 P
                 , 
                 
                 7548
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000001; B = 7'b0010011; // Expected: {'P': 19}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000001; B = 7'b0010011; | Outputs: P=%b | Expected: P=%d",
                 1553,
                 
                 P
                 , 
                 
                 19
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101101; B = 7'b1001100; // Expected: {'P': 8284}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101101; B = 7'b1001100; | Outputs: P=%b | Expected: P=%d",
                 1554,
                 
                 P
                 , 
                 
                 8284
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101010; B = 7'b1011100; // Expected: {'P': 3864}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101010; B = 7'b1011100; | Outputs: P=%b | Expected: P=%d",
                 1555,
                 
                 P
                 , 
                 
                 3864
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010001; B = 7'b0001100; // Expected: {'P': 972}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010001; B = 7'b0001100; | Outputs: P=%b | Expected: P=%d",
                 1556,
                 
                 P
                 , 
                 
                 972
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100110; B = 7'b1010110; // Expected: {'P': 8772}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100110; B = 7'b1010110; | Outputs: P=%b | Expected: P=%d",
                 1557,
                 
                 P
                 , 
                 
                 8772
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001100; B = 7'b0100101; // Expected: {'P': 444}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001100; B = 7'b0100101; | Outputs: P=%b | Expected: P=%d",
                 1558,
                 
                 P
                 , 
                 
                 444
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011000; B = 7'b1011101; // Expected: {'P': 2232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011000; B = 7'b1011101; | Outputs: P=%b | Expected: P=%d",
                 1559,
                 
                 P
                 , 
                 
                 2232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111000; B = 7'b1101101; // Expected: {'P': 13080}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111000; B = 7'b1101101; | Outputs: P=%b | Expected: P=%d",
                 1560,
                 
                 P
                 , 
                 
                 13080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000000; B = 7'b0010100; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000000; B = 7'b0010100; | Outputs: P=%b | Expected: P=%d",
                 1561,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000110; B = 7'b0000101; // Expected: {'P': 350}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000110; B = 7'b0000101; | Outputs: P=%b | Expected: P=%d",
                 1562,
                 
                 P
                 , 
                 
                 350
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111000; B = 7'b0101011; // Expected: {'P': 5160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111000; B = 7'b0101011; | Outputs: P=%b | Expected: P=%d",
                 1563,
                 
                 P
                 , 
                 
                 5160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100110; B = 7'b1011001; // Expected: {'P': 9078}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100110; B = 7'b1011001; | Outputs: P=%b | Expected: P=%d",
                 1564,
                 
                 P
                 , 
                 
                 9078
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101111; B = 7'b1000110; // Expected: {'P': 3290}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101111; B = 7'b1000110; | Outputs: P=%b | Expected: P=%d",
                 1565,
                 
                 P
                 , 
                 
                 3290
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010000; B = 7'b0111001; // Expected: {'P': 912}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010000; B = 7'b0111001; | Outputs: P=%b | Expected: P=%d",
                 1566,
                 
                 P
                 , 
                 
                 912
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111000; B = 7'b1010010; // Expected: {'P': 9840}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111000; B = 7'b1010010; | Outputs: P=%b | Expected: P=%d",
                 1567,
                 
                 P
                 , 
                 
                 9840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110100; B = 7'b0100011; // Expected: {'P': 4060}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110100; B = 7'b0100011; | Outputs: P=%b | Expected: P=%d",
                 1568,
                 
                 P
                 , 
                 
                 4060
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000101; B = 7'b1111100; // Expected: {'P': 8556}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000101; B = 7'b1111100; | Outputs: P=%b | Expected: P=%d",
                 1569,
                 
                 P
                 , 
                 
                 8556
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001001; B = 7'b1010100; // Expected: {'P': 756}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001001; B = 7'b1010100; | Outputs: P=%b | Expected: P=%d",
                 1570,
                 
                 P
                 , 
                 
                 756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110101; B = 7'b1001111; // Expected: {'P': 9243}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110101; B = 7'b1001111; | Outputs: P=%b | Expected: P=%d",
                 1571,
                 
                 P
                 , 
                 
                 9243
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111001; B = 7'b0101100; // Expected: {'P': 5324}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111001; B = 7'b0101100; | Outputs: P=%b | Expected: P=%d",
                 1572,
                 
                 P
                 , 
                 
                 5324
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101101; B = 7'b1111101; // Expected: {'P': 13625}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101101; B = 7'b1111101; | Outputs: P=%b | Expected: P=%d",
                 1573,
                 
                 P
                 , 
                 
                 13625
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111001; B = 7'b0101101; // Expected: {'P': 5445}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111001; B = 7'b0101101; | Outputs: P=%b | Expected: P=%d",
                 1574,
                 
                 P
                 , 
                 
                 5445
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010110; B = 7'b1011001; // Expected: {'P': 7654}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010110; B = 7'b1011001; | Outputs: P=%b | Expected: P=%d",
                 1575,
                 
                 P
                 , 
                 
                 7654
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101101; B = 7'b0001001; // Expected: {'P': 405}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101101; B = 7'b0001001; | Outputs: P=%b | Expected: P=%d",
                 1576,
                 
                 P
                 , 
                 
                 405
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011001; B = 7'b0011010; // Expected: {'P': 650}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011001; B = 7'b0011010; | Outputs: P=%b | Expected: P=%d",
                 1577,
                 
                 P
                 , 
                 
                 650
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110100; B = 7'b1010010; // Expected: {'P': 9512}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110100; B = 7'b1010010; | Outputs: P=%b | Expected: P=%d",
                 1578,
                 
                 P
                 , 
                 
                 9512
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110000; B = 7'b1011101; // Expected: {'P': 4464}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110000; B = 7'b1011101; | Outputs: P=%b | Expected: P=%d",
                 1579,
                 
                 P
                 , 
                 
                 4464
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001000; B = 7'b1001111; // Expected: {'P': 5688}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001000; B = 7'b1001111; | Outputs: P=%b | Expected: P=%d",
                 1580,
                 
                 P
                 , 
                 
                 5688
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101101; B = 7'b0001001; // Expected: {'P': 981}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101101; B = 7'b0001001; | Outputs: P=%b | Expected: P=%d",
                 1581,
                 
                 P
                 , 
                 
                 981
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110010; B = 7'b1100001; // Expected: {'P': 11058}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110010; B = 7'b1100001; | Outputs: P=%b | Expected: P=%d",
                 1582,
                 
                 P
                 , 
                 
                 11058
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110100; B = 7'b1010100; // Expected: {'P': 9744}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110100; B = 7'b1010100; | Outputs: P=%b | Expected: P=%d",
                 1583,
                 
                 P
                 , 
                 
                 9744
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011001; B = 7'b1001011; // Expected: {'P': 6675}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011001; B = 7'b1001011; | Outputs: P=%b | Expected: P=%d",
                 1584,
                 
                 P
                 , 
                 
                 6675
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000001; B = 7'b1011010; // Expected: {'P': 90}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000001; B = 7'b1011010; | Outputs: P=%b | Expected: P=%d",
                 1585,
                 
                 P
                 , 
                 
                 90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001110; B = 7'b1110111; // Expected: {'P': 1666}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001110; B = 7'b1110111; | Outputs: P=%b | Expected: P=%d",
                 1586,
                 
                 P
                 , 
                 
                 1666
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001110; B = 7'b0101110; // Expected: {'P': 3588}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001110; B = 7'b0101110; | Outputs: P=%b | Expected: P=%d",
                 1587,
                 
                 P
                 , 
                 
                 3588
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000011; B = 7'b1001001; // Expected: {'P': 219}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000011; B = 7'b1001001; | Outputs: P=%b | Expected: P=%d",
                 1588,
                 
                 P
                 , 
                 
                 219
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010110; B = 7'b0001000; // Expected: {'P': 176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010110; B = 7'b0001000; | Outputs: P=%b | Expected: P=%d",
                 1589,
                 
                 P
                 , 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000110; B = 7'b1010111; // Expected: {'P': 6090}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000110; B = 7'b1010111; | Outputs: P=%b | Expected: P=%d",
                 1590,
                 
                 P
                 , 
                 
                 6090
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000101; B = 7'b0110011; // Expected: {'P': 3519}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000101; B = 7'b0110011; | Outputs: P=%b | Expected: P=%d",
                 1591,
                 
                 P
                 , 
                 
                 3519
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001100; B = 7'b1000110; // Expected: {'P': 840}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001100; B = 7'b1000110; | Outputs: P=%b | Expected: P=%d",
                 1592,
                 
                 P
                 , 
                 
                 840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111110; B = 7'b0110011; // Expected: {'P': 3162}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111110; B = 7'b0110011; | Outputs: P=%b | Expected: P=%d",
                 1593,
                 
                 P
                 , 
                 
                 3162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111000; B = 7'b1011000; // Expected: {'P': 4928}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111000; B = 7'b1011000; | Outputs: P=%b | Expected: P=%d",
                 1594,
                 
                 P
                 , 
                 
                 4928
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010010; B = 7'b1000000; // Expected: {'P': 5248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010010; B = 7'b1000000; | Outputs: P=%b | Expected: P=%d",
                 1595,
                 
                 P
                 , 
                 
                 5248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101110; B = 7'b1001000; // Expected: {'P': 7920}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101110; B = 7'b1001000; | Outputs: P=%b | Expected: P=%d",
                 1596,
                 
                 P
                 , 
                 
                 7920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000110; B = 7'b0010100; // Expected: {'P': 120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000110; B = 7'b0010100; | Outputs: P=%b | Expected: P=%d",
                 1597,
                 
                 P
                 , 
                 
                 120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101111; B = 7'b1111100; // Expected: {'P': 13764}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101111; B = 7'b1111100; | Outputs: P=%b | Expected: P=%d",
                 1598,
                 
                 P
                 , 
                 
                 13764
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101111; B = 7'b1001110; // Expected: {'P': 3666}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101111; B = 7'b1001110; | Outputs: P=%b | Expected: P=%d",
                 1599,
                 
                 P
                 , 
                 
                 3666
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010101; B = 7'b1001111; // Expected: {'P': 6715}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010101; B = 7'b1001111; | Outputs: P=%b | Expected: P=%d",
                 1600,
                 
                 P
                 , 
                 
                 6715
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000111; B = 7'b1001010; // Expected: {'P': 518}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000111; B = 7'b1001010; | Outputs: P=%b | Expected: P=%d",
                 1601,
                 
                 P
                 , 
                 
                 518
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111010; B = 7'b0001000; // Expected: {'P': 976}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111010; B = 7'b0001000; | Outputs: P=%b | Expected: P=%d",
                 1602,
                 
                 P
                 , 
                 
                 976
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101100; B = 7'b0011011; // Expected: {'P': 2916}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101100; B = 7'b0011011; | Outputs: P=%b | Expected: P=%d",
                 1603,
                 
                 P
                 , 
                 
                 2916
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001111; B = 7'b1000101; // Expected: {'P': 1035}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001111; B = 7'b1000101; | Outputs: P=%b | Expected: P=%d",
                 1604,
                 
                 P
                 , 
                 
                 1035
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011100; B = 7'b0000100; // Expected: {'P': 368}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011100; B = 7'b0000100; | Outputs: P=%b | Expected: P=%d",
                 1605,
                 
                 P
                 , 
                 
                 368
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110111; B = 7'b0010000; // Expected: {'P': 880}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110111; B = 7'b0010000; | Outputs: P=%b | Expected: P=%d",
                 1606,
                 
                 P
                 , 
                 
                 880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101110; B = 7'b0100110; // Expected: {'P': 1748}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101110; B = 7'b0100110; | Outputs: P=%b | Expected: P=%d",
                 1607,
                 
                 P
                 , 
                 
                 1748
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000000; B = 7'b1111101; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000000; B = 7'b1111101; | Outputs: P=%b | Expected: P=%d",
                 1608,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000011; B = 7'b1100111; // Expected: {'P': 6901}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000011; B = 7'b1100111; | Outputs: P=%b | Expected: P=%d",
                 1609,
                 
                 P
                 , 
                 
                 6901
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001111; B = 7'b0011101; // Expected: {'P': 2291}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001111; B = 7'b0011101; | Outputs: P=%b | Expected: P=%d",
                 1610,
                 
                 P
                 , 
                 
                 2291
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001101; B = 7'b0010000; // Expected: {'P': 1232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001101; B = 7'b0010000; | Outputs: P=%b | Expected: P=%d",
                 1611,
                 
                 P
                 , 
                 
                 1232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110100; B = 7'b0011100; // Expected: {'P': 1456}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110100; B = 7'b0011100; | Outputs: P=%b | Expected: P=%d",
                 1612,
                 
                 P
                 , 
                 
                 1456
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100100; B = 7'b1010111; // Expected: {'P': 3132}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100100; B = 7'b1010111; | Outputs: P=%b | Expected: P=%d",
                 1613,
                 
                 P
                 , 
                 
                 3132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000010; B = 7'b1111011; // Expected: {'P': 246}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000010; B = 7'b1111011; | Outputs: P=%b | Expected: P=%d",
                 1614,
                 
                 P
                 , 
                 
                 246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101001; B = 7'b1111001; // Expected: {'P': 12705}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101001; B = 7'b1111001; | Outputs: P=%b | Expected: P=%d",
                 1615,
                 
                 P
                 , 
                 
                 12705
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100110; B = 7'b0110110; // Expected: {'P': 2052}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100110; B = 7'b0110110; | Outputs: P=%b | Expected: P=%d",
                 1616,
                 
                 P
                 , 
                 
                 2052
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110101; B = 7'b0111110; // Expected: {'P': 3286}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110101; B = 7'b0111110; | Outputs: P=%b | Expected: P=%d",
                 1617,
                 
                 P
                 , 
                 
                 3286
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101111; B = 7'b0110010; // Expected: {'P': 5550}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101111; B = 7'b0110010; | Outputs: P=%b | Expected: P=%d",
                 1618,
                 
                 P
                 , 
                 
                 5550
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011101; B = 7'b0001011; // Expected: {'P': 319}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011101; B = 7'b0001011; | Outputs: P=%b | Expected: P=%d",
                 1619,
                 
                 P
                 , 
                 
                 319
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001000; B = 7'b0000110; // Expected: {'P': 48}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001000; B = 7'b0000110; | Outputs: P=%b | Expected: P=%d",
                 1620,
                 
                 P
                 , 
                 
                 48
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111010; B = 7'b0010100; // Expected: {'P': 1160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111010; B = 7'b0010100; | Outputs: P=%b | Expected: P=%d",
                 1621,
                 
                 P
                 , 
                 
                 1160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010100; B = 7'b1100110; // Expected: {'P': 2040}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010100; B = 7'b1100110; | Outputs: P=%b | Expected: P=%d",
                 1622,
                 
                 P
                 , 
                 
                 2040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011100; B = 7'b0101001; // Expected: {'P': 3772}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011100; B = 7'b0101001; | Outputs: P=%b | Expected: P=%d",
                 1623,
                 
                 P
                 , 
                 
                 3772
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011010; B = 7'b1110111; // Expected: {'P': 10710}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011010; B = 7'b1110111; | Outputs: P=%b | Expected: P=%d",
                 1624,
                 
                 P
                 , 
                 
                 10710
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111001; B = 7'b0000110; // Expected: {'P': 726}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111001; B = 7'b0000110; | Outputs: P=%b | Expected: P=%d",
                 1625,
                 
                 P
                 , 
                 
                 726
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100110; B = 7'b1010001; // Expected: {'P': 8262}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100110; B = 7'b1010001; | Outputs: P=%b | Expected: P=%d",
                 1626,
                 
                 P
                 , 
                 
                 8262
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100011; B = 7'b1011010; // Expected: {'P': 3150}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100011; B = 7'b1011010; | Outputs: P=%b | Expected: P=%d",
                 1627,
                 
                 P
                 , 
                 
                 3150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111101; B = 7'b0101011; // Expected: {'P': 2623}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111101; B = 7'b0101011; | Outputs: P=%b | Expected: P=%d",
                 1628,
                 
                 P
                 , 
                 
                 2623
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010001; B = 7'b0101101; // Expected: {'P': 765}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010001; B = 7'b0101101; | Outputs: P=%b | Expected: P=%d",
                 1629,
                 
                 P
                 , 
                 
                 765
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111101; B = 7'b1001110; // Expected: {'P': 4758}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111101; B = 7'b1001110; | Outputs: P=%b | Expected: P=%d",
                 1630,
                 
                 P
                 , 
                 
                 4758
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001100; B = 7'b0001000; // Expected: {'P': 608}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001100; B = 7'b0001000; | Outputs: P=%b | Expected: P=%d",
                 1631,
                 
                 P
                 , 
                 
                 608
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000111; B = 7'b1111110; // Expected: {'P': 882}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000111; B = 7'b1111110; | Outputs: P=%b | Expected: P=%d",
                 1632,
                 
                 P
                 , 
                 
                 882
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011001; B = 7'b1011100; // Expected: {'P': 8188}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011001; B = 7'b1011100; | Outputs: P=%b | Expected: P=%d",
                 1633,
                 
                 P
                 , 
                 
                 8188
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100110; B = 7'b1010100; // Expected: {'P': 8568}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100110; B = 7'b1010100; | Outputs: P=%b | Expected: P=%d",
                 1634,
                 
                 P
                 , 
                 
                 8568
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110101; B = 7'b0000011; // Expected: {'P': 159}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110101; B = 7'b0000011; | Outputs: P=%b | Expected: P=%d",
                 1635,
                 
                 P
                 , 
                 
                 159
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001000; B = 7'b1010001; // Expected: {'P': 5832}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001000; B = 7'b1010001; | Outputs: P=%b | Expected: P=%d",
                 1636,
                 
                 P
                 , 
                 
                 5832
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010111; B = 7'b1010000; // Expected: {'P': 1840}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010111; B = 7'b1010000; | Outputs: P=%b | Expected: P=%d",
                 1637,
                 
                 P
                 , 
                 
                 1840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101101; B = 7'b1111011; // Expected: {'P': 13407}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101101; B = 7'b1111011; | Outputs: P=%b | Expected: P=%d",
                 1638,
                 
                 P
                 , 
                 
                 13407
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011010; B = 7'b0000101; // Expected: {'P': 450}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011010; B = 7'b0000101; | Outputs: P=%b | Expected: P=%d",
                 1639,
                 
                 P
                 , 
                 
                 450
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000101; B = 7'b1100011; // Expected: {'P': 6831}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000101; B = 7'b1100011; | Outputs: P=%b | Expected: P=%d",
                 1640,
                 
                 P
                 , 
                 
                 6831
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110100; B = 7'b0100100; // Expected: {'P': 1872}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110100; B = 7'b0100100; | Outputs: P=%b | Expected: P=%d",
                 1641,
                 
                 P
                 , 
                 
                 1872
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101110; B = 7'b0000001; // Expected: {'P': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101110; B = 7'b0000001; | Outputs: P=%b | Expected: P=%d",
                 1642,
                 
                 P
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101110; B = 7'b1001011; // Expected: {'P': 3450}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101110; B = 7'b1001011; | Outputs: P=%b | Expected: P=%d",
                 1643,
                 
                 P
                 , 
                 
                 3450
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010000; B = 7'b0100111; // Expected: {'P': 624}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010000; B = 7'b0100111; | Outputs: P=%b | Expected: P=%d",
                 1644,
                 
                 P
                 , 
                 
                 624
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101011; B = 7'b1110101; // Expected: {'P': 5031}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101011; B = 7'b1110101; | Outputs: P=%b | Expected: P=%d",
                 1645,
                 
                 P
                 , 
                 
                 5031
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100100; B = 7'b1001101; // Expected: {'P': 2772}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100100; B = 7'b1001101; | Outputs: P=%b | Expected: P=%d",
                 1646,
                 
                 P
                 , 
                 
                 2772
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100000; B = 7'b1011001; // Expected: {'P': 8544}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100000; B = 7'b1011001; | Outputs: P=%b | Expected: P=%d",
                 1647,
                 
                 P
                 , 
                 
                 8544
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100111; B = 7'b1110001; // Expected: {'P': 4407}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100111; B = 7'b1110001; | Outputs: P=%b | Expected: P=%d",
                 1648,
                 
                 P
                 , 
                 
                 4407
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111100; B = 7'b1010000; // Expected: {'P': 4800}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111100; B = 7'b1010000; | Outputs: P=%b | Expected: P=%d",
                 1649,
                 
                 P
                 , 
                 
                 4800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010100; B = 7'b1001111; // Expected: {'P': 1580}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010100; B = 7'b1001111; | Outputs: P=%b | Expected: P=%d",
                 1650,
                 
                 P
                 , 
                 
                 1580
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001000; B = 7'b1101011; // Expected: {'P': 856}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001000; B = 7'b1101011; | Outputs: P=%b | Expected: P=%d",
                 1651,
                 
                 P
                 , 
                 
                 856
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110111; B = 7'b1100011; // Expected: {'P': 11781}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110111; B = 7'b1100011; | Outputs: P=%b | Expected: P=%d",
                 1652,
                 
                 P
                 , 
                 
                 11781
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001001; B = 7'b1001000; // Expected: {'P': 5256}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001001; B = 7'b1001000; | Outputs: P=%b | Expected: P=%d",
                 1653,
                 
                 P
                 , 
                 
                 5256
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110001; B = 7'b0010101; // Expected: {'P': 1029}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110001; B = 7'b0010101; | Outputs: P=%b | Expected: P=%d",
                 1654,
                 
                 P
                 , 
                 
                 1029
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110100; B = 7'b1100111; // Expected: {'P': 5356}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110100; B = 7'b1100111; | Outputs: P=%b | Expected: P=%d",
                 1655,
                 
                 P
                 , 
                 
                 5356
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011100; B = 7'b0010100; // Expected: {'P': 1840}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011100; B = 7'b0010100; | Outputs: P=%b | Expected: P=%d",
                 1656,
                 
                 P
                 , 
                 
                 1840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010010; B = 7'b1110010; // Expected: {'P': 2052}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010010; B = 7'b1110010; | Outputs: P=%b | Expected: P=%d",
                 1657,
                 
                 P
                 , 
                 
                 2052
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010010; B = 7'b1100111; // Expected: {'P': 1854}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010010; B = 7'b1100111; | Outputs: P=%b | Expected: P=%d",
                 1658,
                 
                 P
                 , 
                 
                 1854
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001000; B = 7'b1100101; // Expected: {'P': 808}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001000; B = 7'b1100101; | Outputs: P=%b | Expected: P=%d",
                 1659,
                 
                 P
                 , 
                 
                 808
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011100; B = 7'b1100011; // Expected: {'P': 2772}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011100; B = 7'b1100011; | Outputs: P=%b | Expected: P=%d",
                 1660,
                 
                 P
                 , 
                 
                 2772
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101010; B = 7'b1101101; // Expected: {'P': 4578}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101010; B = 7'b1101101; | Outputs: P=%b | Expected: P=%d",
                 1661,
                 
                 P
                 , 
                 
                 4578
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011101; B = 7'b0011000; // Expected: {'P': 696}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011101; B = 7'b0011000; | Outputs: P=%b | Expected: P=%d",
                 1662,
                 
                 P
                 , 
                 
                 696
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100111; B = 7'b0100010; // Expected: {'P': 1326}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100111; B = 7'b0100010; | Outputs: P=%b | Expected: P=%d",
                 1663,
                 
                 P
                 , 
                 
                 1326
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110010; B = 7'b0111111; // Expected: {'P': 3150}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110010; B = 7'b0111111; | Outputs: P=%b | Expected: P=%d",
                 1664,
                 
                 P
                 , 
                 
                 3150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111100; B = 7'b1001101; // Expected: {'P': 4620}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111100; B = 7'b1001101; | Outputs: P=%b | Expected: P=%d",
                 1665,
                 
                 P
                 , 
                 
                 4620
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000010; B = 7'b0010011; // Expected: {'P': 1254}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000010; B = 7'b0010011; | Outputs: P=%b | Expected: P=%d",
                 1666,
                 
                 P
                 , 
                 
                 1254
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001110; B = 7'b1111100; // Expected: {'P': 9672}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001110; B = 7'b1111100; | Outputs: P=%b | Expected: P=%d",
                 1667,
                 
                 P
                 , 
                 
                 9672
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011101; B = 7'b1110110; // Expected: {'P': 3422}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011101; B = 7'b1110110; | Outputs: P=%b | Expected: P=%d",
                 1668,
                 
                 P
                 , 
                 
                 3422
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001001; B = 7'b1000110; // Expected: {'P': 5110}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001001; B = 7'b1000110; | Outputs: P=%b | Expected: P=%d",
                 1669,
                 
                 P
                 , 
                 
                 5110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110000; B = 7'b0110011; // Expected: {'P': 2448}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110000; B = 7'b0110011; | Outputs: P=%b | Expected: P=%d",
                 1670,
                 
                 P
                 , 
                 
                 2448
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111100; B = 7'b1101111; // Expected: {'P': 6660}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111100; B = 7'b1101111; | Outputs: P=%b | Expected: P=%d",
                 1671,
                 
                 P
                 , 
                 
                 6660
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011011; B = 7'b1000100; // Expected: {'P': 6188}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011011; B = 7'b1000100; | Outputs: P=%b | Expected: P=%d",
                 1672,
                 
                 P
                 , 
                 
                 6188
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101100; B = 7'b1110111; // Expected: {'P': 12852}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101100; B = 7'b1110111; | Outputs: P=%b | Expected: P=%d",
                 1673,
                 
                 P
                 , 
                 
                 12852
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101011; B = 7'b0010001; // Expected: {'P': 731}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101011; B = 7'b0010001; | Outputs: P=%b | Expected: P=%d",
                 1674,
                 
                 P
                 , 
                 
                 731
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011010; B = 7'b1100000; // Expected: {'P': 2496}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011010; B = 7'b1100000; | Outputs: P=%b | Expected: P=%d",
                 1675,
                 
                 P
                 , 
                 
                 2496
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110110; B = 7'b0100010; // Expected: {'P': 1836}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110110; B = 7'b0100010; | Outputs: P=%b | Expected: P=%d",
                 1676,
                 
                 P
                 , 
                 
                 1836
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101000; B = 7'b0100111; // Expected: {'P': 4056}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101000; B = 7'b0100111; | Outputs: P=%b | Expected: P=%d",
                 1677,
                 
                 P
                 , 
                 
                 4056
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011010; B = 7'b0111100; // Expected: {'P': 1560}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011010; B = 7'b0111100; | Outputs: P=%b | Expected: P=%d",
                 1678,
                 
                 P
                 , 
                 
                 1560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111001; B = 7'b1101001; // Expected: {'P': 5985}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111001; B = 7'b1101001; | Outputs: P=%b | Expected: P=%d",
                 1679,
                 
                 P
                 , 
                 
                 5985
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011010; B = 7'b1000000; // Expected: {'P': 1664}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011010; B = 7'b1000000; | Outputs: P=%b | Expected: P=%d",
                 1680,
                 
                 P
                 , 
                 
                 1664
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101011; B = 7'b1011010; // Expected: {'P': 9630}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101011; B = 7'b1011010; | Outputs: P=%b | Expected: P=%d",
                 1681,
                 
                 P
                 , 
                 
                 9630
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010011; B = 7'b1011101; // Expected: {'P': 1767}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010011; B = 7'b1011101; | Outputs: P=%b | Expected: P=%d",
                 1682,
                 
                 P
                 , 
                 
                 1767
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000111; B = 7'b1101100; // Expected: {'P': 756}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000111; B = 7'b1101100; | Outputs: P=%b | Expected: P=%d",
                 1683,
                 
                 P
                 , 
                 
                 756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110100; B = 7'b1001010; // Expected: {'P': 3848}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110100; B = 7'b1001010; | Outputs: P=%b | Expected: P=%d",
                 1684,
                 
                 P
                 , 
                 
                 3848
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111100; B = 7'b0111111; // Expected: {'P': 3780}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111100; B = 7'b0111111; | Outputs: P=%b | Expected: P=%d",
                 1685,
                 
                 P
                 , 
                 
                 3780
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001001; B = 7'b1001010; // Expected: {'P': 5402}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001001; B = 7'b1001010; | Outputs: P=%b | Expected: P=%d",
                 1686,
                 
                 P
                 , 
                 
                 5402
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100010; B = 7'b1001101; // Expected: {'P': 2618}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100010; B = 7'b1001101; | Outputs: P=%b | Expected: P=%d",
                 1687,
                 
                 P
                 , 
                 
                 2618
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111100; B = 7'b1001010; // Expected: {'P': 4440}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111100; B = 7'b1001010; | Outputs: P=%b | Expected: P=%d",
                 1688,
                 
                 P
                 , 
                 
                 4440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111110; B = 7'b1111101; // Expected: {'P': 15750}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111110; B = 7'b1111101; | Outputs: P=%b | Expected: P=%d",
                 1689,
                 
                 P
                 , 
                 
                 15750
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100010; B = 7'b0000101; // Expected: {'P': 490}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100010; B = 7'b0000101; | Outputs: P=%b | Expected: P=%d",
                 1690,
                 
                 P
                 , 
                 
                 490
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011001; B = 7'b1001101; // Expected: {'P': 6853}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011001; B = 7'b1001101; | Outputs: P=%b | Expected: P=%d",
                 1691,
                 
                 P
                 , 
                 
                 6853
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010000; B = 7'b0011010; // Expected: {'P': 2080}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010000; B = 7'b0011010; | Outputs: P=%b | Expected: P=%d",
                 1692,
                 
                 P
                 , 
                 
                 2080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000100; B = 7'b0100100; // Expected: {'P': 144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000100; B = 7'b0100100; | Outputs: P=%b | Expected: P=%d",
                 1693,
                 
                 P
                 , 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001110; B = 7'b0000111; // Expected: {'P': 546}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001110; B = 7'b0000111; | Outputs: P=%b | Expected: P=%d",
                 1694,
                 
                 P
                 , 
                 
                 546
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001011; B = 7'b0010111; // Expected: {'P': 253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001011; B = 7'b0010111; | Outputs: P=%b | Expected: P=%d",
                 1695,
                 
                 P
                 , 
                 
                 253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101010; B = 7'b1101110; // Expected: {'P': 4620}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101010; B = 7'b1101110; | Outputs: P=%b | Expected: P=%d",
                 1696,
                 
                 P
                 , 
                 
                 4620
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101011; B = 7'b1010110; // Expected: {'P': 3698}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101011; B = 7'b1010110; | Outputs: P=%b | Expected: P=%d",
                 1697,
                 
                 P
                 , 
                 
                 3698
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111100; B = 7'b1011001; // Expected: {'P': 11036}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111100; B = 7'b1011001; | Outputs: P=%b | Expected: P=%d",
                 1698,
                 
                 P
                 , 
                 
                 11036
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011101; B = 7'b0000010; // Expected: {'P': 58}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011101; B = 7'b0000010; | Outputs: P=%b | Expected: P=%d",
                 1699,
                 
                 P
                 , 
                 
                 58
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110010; B = 7'b1011011; // Expected: {'P': 4550}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110010; B = 7'b1011011; | Outputs: P=%b | Expected: P=%d",
                 1700,
                 
                 P
                 , 
                 
                 4550
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101100; B = 7'b0011101; // Expected: {'P': 3132}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101100; B = 7'b0011101; | Outputs: P=%b | Expected: P=%d",
                 1701,
                 
                 P
                 , 
                 
                 3132
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110111; B = 7'b0100000; // Expected: {'P': 3808}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110111; B = 7'b0100000; | Outputs: P=%b | Expected: P=%d",
                 1702,
                 
                 P
                 , 
                 
                 3808
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111100; B = 7'b0101000; // Expected: {'P': 2400}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111100; B = 7'b0101000; | Outputs: P=%b | Expected: P=%d",
                 1703,
                 
                 P
                 , 
                 
                 2400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101000; B = 7'b0110011; // Expected: {'P': 2040}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101000; B = 7'b0110011; | Outputs: P=%b | Expected: P=%d",
                 1704,
                 
                 P
                 , 
                 
                 2040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001011; B = 7'b1111001; // Expected: {'P': 1331}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001011; B = 7'b1111001; | Outputs: P=%b | Expected: P=%d",
                 1705,
                 
                 P
                 , 
                 
                 1331
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110100; B = 7'b1100111; // Expected: {'P': 11948}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110100; B = 7'b1100111; | Outputs: P=%b | Expected: P=%d",
                 1706,
                 
                 P
                 , 
                 
                 11948
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101111; B = 7'b1011110; // Expected: {'P': 4418}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101111; B = 7'b1011110; | Outputs: P=%b | Expected: P=%d",
                 1707,
                 
                 P
                 , 
                 
                 4418
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110000; B = 7'b1000010; // Expected: {'P': 7392}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110000; B = 7'b1000010; | Outputs: P=%b | Expected: P=%d",
                 1708,
                 
                 P
                 , 
                 
                 7392
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101100; B = 7'b0101000; // Expected: {'P': 4320}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101100; B = 7'b0101000; | Outputs: P=%b | Expected: P=%d",
                 1709,
                 
                 P
                 , 
                 
                 4320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001010; B = 7'b0011100; // Expected: {'P': 2072}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001010; B = 7'b0011100; | Outputs: P=%b | Expected: P=%d",
                 1710,
                 
                 P
                 , 
                 
                 2072
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000101; B = 7'b0111001; // Expected: {'P': 3933}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000101; B = 7'b0111001; | Outputs: P=%b | Expected: P=%d",
                 1711,
                 
                 P
                 , 
                 
                 3933
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100001; B = 7'b1010111; // Expected: {'P': 8439}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100001; B = 7'b1010111; | Outputs: P=%b | Expected: P=%d",
                 1712,
                 
                 P
                 , 
                 
                 8439
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000011; B = 7'b1000001; // Expected: {'P': 4355}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000011; B = 7'b1000001; | Outputs: P=%b | Expected: P=%d",
                 1713,
                 
                 P
                 , 
                 
                 4355
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111101; B = 7'b0001111; // Expected: {'P': 915}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111101; B = 7'b0001111; | Outputs: P=%b | Expected: P=%d",
                 1714,
                 
                 P
                 , 
                 
                 915
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011011; B = 7'b0111110; // Expected: {'P': 1674}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011011; B = 7'b0111110; | Outputs: P=%b | Expected: P=%d",
                 1715,
                 
                 P
                 , 
                 
                 1674
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100001; B = 7'b0010100; // Expected: {'P': 660}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100001; B = 7'b0010100; | Outputs: P=%b | Expected: P=%d",
                 1716,
                 
                 P
                 , 
                 
                 660
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000010; B = 7'b0000110; // Expected: {'P': 12}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000010; B = 7'b0000110; | Outputs: P=%b | Expected: P=%d",
                 1717,
                 
                 P
                 , 
                 
                 12
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111000; B = 7'b1111000; // Expected: {'P': 6720}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111000; B = 7'b1111000; | Outputs: P=%b | Expected: P=%d",
                 1718,
                 
                 P
                 , 
                 
                 6720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000110; B = 7'b1010000; // Expected: {'P': 5600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000110; B = 7'b1010000; | Outputs: P=%b | Expected: P=%d",
                 1719,
                 
                 P
                 , 
                 
                 5600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110011; B = 7'b0011111; // Expected: {'P': 1581}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110011; B = 7'b0011111; | Outputs: P=%b | Expected: P=%d",
                 1720,
                 
                 P
                 , 
                 
                 1581
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110101; B = 7'b0011010; // Expected: {'P': 3042}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110101; B = 7'b0011010; | Outputs: P=%b | Expected: P=%d",
                 1721,
                 
                 P
                 , 
                 
                 3042
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101100; B = 7'b0111111; // Expected: {'P': 6804}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101100; B = 7'b0111111; | Outputs: P=%b | Expected: P=%d",
                 1722,
                 
                 P
                 , 
                 
                 6804
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000101; B = 7'b0111100; // Expected: {'P': 300}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000101; B = 7'b0111100; | Outputs: P=%b | Expected: P=%d",
                 1723,
                 
                 P
                 , 
                 
                 300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010000; B = 7'b1101000; // Expected: {'P': 1664}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010000; B = 7'b1101000; | Outputs: P=%b | Expected: P=%d",
                 1724,
                 
                 P
                 , 
                 
                 1664
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101101; B = 7'b0111100; // Expected: {'P': 6540}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101101; B = 7'b0111100; | Outputs: P=%b | Expected: P=%d",
                 1725,
                 
                 P
                 , 
                 
                 6540
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011101; B = 7'b0100011; // Expected: {'P': 1015}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011101; B = 7'b0100011; | Outputs: P=%b | Expected: P=%d",
                 1726,
                 
                 P
                 , 
                 
                 1015
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111111; B = 7'b0110011; // Expected: {'P': 3213}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111111; B = 7'b0110011; | Outputs: P=%b | Expected: P=%d",
                 1727,
                 
                 P
                 , 
                 
                 3213
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110100; B = 7'b1001100; // Expected: {'P': 8816}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110100; B = 7'b1001100; | Outputs: P=%b | Expected: P=%d",
                 1728,
                 
                 P
                 , 
                 
                 8816
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000101; B = 7'b0101110; // Expected: {'P': 3174}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000101; B = 7'b0101110; | Outputs: P=%b | Expected: P=%d",
                 1729,
                 
                 P
                 , 
                 
                 3174
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010000; B = 7'b1000110; // Expected: {'P': 5600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010000; B = 7'b1000110; | Outputs: P=%b | Expected: P=%d",
                 1730,
                 
                 P
                 , 
                 
                 5600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010111; B = 7'b0001011; // Expected: {'P': 957}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010111; B = 7'b0001011; | Outputs: P=%b | Expected: P=%d",
                 1731,
                 
                 P
                 , 
                 
                 957
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010101; B = 7'b1110111; // Expected: {'P': 2499}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010101; B = 7'b1110111; | Outputs: P=%b | Expected: P=%d",
                 1732,
                 
                 P
                 , 
                 
                 2499
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111000; B = 7'b1101001; // Expected: {'P': 12600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111000; B = 7'b1101001; | Outputs: P=%b | Expected: P=%d",
                 1733,
                 
                 P
                 , 
                 
                 12600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010011; B = 7'b0100000; // Expected: {'P': 2656}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010011; B = 7'b0100000; | Outputs: P=%b | Expected: P=%d",
                 1734,
                 
                 P
                 , 
                 
                 2656
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101011; B = 7'b0010100; // Expected: {'P': 2140}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101011; B = 7'b0010100; | Outputs: P=%b | Expected: P=%d",
                 1735,
                 
                 P
                 , 
                 
                 2140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111000; B = 7'b0000101; // Expected: {'P': 600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111000; B = 7'b0000101; | Outputs: P=%b | Expected: P=%d",
                 1736,
                 
                 P
                 , 
                 
                 600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110110; B = 7'b0101000; // Expected: {'P': 2160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110110; B = 7'b0101000; | Outputs: P=%b | Expected: P=%d",
                 1737,
                 
                 P
                 , 
                 
                 2160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110011; B = 7'b1100011; // Expected: {'P': 5049}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110011; B = 7'b1100011; | Outputs: P=%b | Expected: P=%d",
                 1738,
                 
                 P
                 , 
                 
                 5049
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010101; B = 7'b1001001; // Expected: {'P': 6205}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010101; B = 7'b1001001; | Outputs: P=%b | Expected: P=%d",
                 1739,
                 
                 P
                 , 
                 
                 6205
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100000; B = 7'b1000011; // Expected: {'P': 6432}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100000; B = 7'b1000011; | Outputs: P=%b | Expected: P=%d",
                 1740,
                 
                 P
                 , 
                 
                 6432
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110011; B = 7'b0011010; // Expected: {'P': 2990}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110011; B = 7'b0011010; | Outputs: P=%b | Expected: P=%d",
                 1741,
                 
                 P
                 , 
                 
                 2990
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111110; B = 7'b1010111; // Expected: {'P': 5394}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111110; B = 7'b1010111; | Outputs: P=%b | Expected: P=%d",
                 1742,
                 
                 P
                 , 
                 
                 5394
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001001; B = 7'b1101011; // Expected: {'P': 963}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001001; B = 7'b1101011; | Outputs: P=%b | Expected: P=%d",
                 1743,
                 
                 P
                 , 
                 
                 963
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011011; B = 7'b1111000; // Expected: {'P': 10920}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011011; B = 7'b1111000; | Outputs: P=%b | Expected: P=%d",
                 1744,
                 
                 P
                 , 
                 
                 10920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011101; B = 7'b0100000; // Expected: {'P': 928}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011101; B = 7'b0100000; | Outputs: P=%b | Expected: P=%d",
                 1745,
                 
                 P
                 , 
                 
                 928
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111111; B = 7'b0000100; // Expected: {'P': 508}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111111; B = 7'b0000100; | Outputs: P=%b | Expected: P=%d",
                 1746,
                 
                 P
                 , 
                 
                 508
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001010; B = 7'b0111110; // Expected: {'P': 4588}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001010; B = 7'b0111110; | Outputs: P=%b | Expected: P=%d",
                 1747,
                 
                 P
                 , 
                 
                 4588
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110101; B = 7'b0100101; // Expected: {'P': 4329}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110101; B = 7'b0100101; | Outputs: P=%b | Expected: P=%d",
                 1748,
                 
                 P
                 , 
                 
                 4329
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001011; B = 7'b0111011; // Expected: {'P': 4425}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001011; B = 7'b0111011; | Outputs: P=%b | Expected: P=%d",
                 1749,
                 
                 P
                 , 
                 
                 4425
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001011; B = 7'b1100110; // Expected: {'P': 1122}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001011; B = 7'b1100110; | Outputs: P=%b | Expected: P=%d",
                 1750,
                 
                 P
                 , 
                 
                 1122
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011101; B = 7'b0100001; // Expected: {'P': 3069}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011101; B = 7'b0100001; | Outputs: P=%b | Expected: P=%d",
                 1751,
                 
                 P
                 , 
                 
                 3069
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100110; B = 7'b0111101; // Expected: {'P': 6222}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100110; B = 7'b0111101; | Outputs: P=%b | Expected: P=%d",
                 1752,
                 
                 P
                 , 
                 
                 6222
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010111; B = 7'b1111000; // Expected: {'P': 2760}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010111; B = 7'b1111000; | Outputs: P=%b | Expected: P=%d",
                 1753,
                 
                 P
                 , 
                 
                 2760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010110; B = 7'b0111100; // Expected: {'P': 5160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010110; B = 7'b0111100; | Outputs: P=%b | Expected: P=%d",
                 1754,
                 
                 P
                 , 
                 
                 5160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110011; B = 7'b0000011; // Expected: {'P': 153}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110011; B = 7'b0000011; | Outputs: P=%b | Expected: P=%d",
                 1755,
                 
                 P
                 , 
                 
                 153
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111100; B = 7'b0110010; // Expected: {'P': 6200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111100; B = 7'b0110010; | Outputs: P=%b | Expected: P=%d",
                 1756,
                 
                 P
                 , 
                 
                 6200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111100; B = 7'b0001001; // Expected: {'P': 1116}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111100; B = 7'b0001001; | Outputs: P=%b | Expected: P=%d",
                 1757,
                 
                 P
                 , 
                 
                 1116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011110; B = 7'b0011001; // Expected: {'P': 2350}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011110; B = 7'b0011001; | Outputs: P=%b | Expected: P=%d",
                 1758,
                 
                 P
                 , 
                 
                 2350
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000010; B = 7'b1011101; // Expected: {'P': 6138}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000010; B = 7'b1011101; | Outputs: P=%b | Expected: P=%d",
                 1759,
                 
                 P
                 , 
                 
                 6138
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010001; B = 7'b1010100; // Expected: {'P': 1428}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010001; B = 7'b1010100; | Outputs: P=%b | Expected: P=%d",
                 1760,
                 
                 P
                 , 
                 
                 1428
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111001; B = 7'b1110010; // Expected: {'P': 6498}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111001; B = 7'b1110010; | Outputs: P=%b | Expected: P=%d",
                 1761,
                 
                 P
                 , 
                 
                 6498
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011101; B = 7'b1010000; // Expected: {'P': 7440}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011101; B = 7'b1010000; | Outputs: P=%b | Expected: P=%d",
                 1762,
                 
                 P
                 , 
                 
                 7440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010101; B = 7'b1100101; // Expected: {'P': 8585}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010101; B = 7'b1100101; | Outputs: P=%b | Expected: P=%d",
                 1763,
                 
                 P
                 , 
                 
                 8585
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110100; B = 7'b0111000; // Expected: {'P': 6496}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110100; B = 7'b0111000; | Outputs: P=%b | Expected: P=%d",
                 1764,
                 
                 P
                 , 
                 
                 6496
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101001; B = 7'b1101010; // Expected: {'P': 4346}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101001; B = 7'b1101010; | Outputs: P=%b | Expected: P=%d",
                 1765,
                 
                 P
                 , 
                 
                 4346
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000110; B = 7'b1011000; // Expected: {'P': 6160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000110; B = 7'b1011000; | Outputs: P=%b | Expected: P=%d",
                 1766,
                 
                 P
                 , 
                 
                 6160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010111; B = 7'b0001001; // Expected: {'P': 207}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010111; B = 7'b0001001; | Outputs: P=%b | Expected: P=%d",
                 1767,
                 
                 P
                 , 
                 
                 207
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010111; B = 7'b0001111; // Expected: {'P': 345}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010111; B = 7'b0001111; | Outputs: P=%b | Expected: P=%d",
                 1768,
                 
                 P
                 , 
                 
                 345
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101111; B = 7'b0001010; // Expected: {'P': 470}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101111; B = 7'b0001010; | Outputs: P=%b | Expected: P=%d",
                 1769,
                 
                 P
                 , 
                 
                 470
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100110; B = 7'b1010010; // Expected: {'P': 8364}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100110; B = 7'b1010010; | Outputs: P=%b | Expected: P=%d",
                 1770,
                 
                 P
                 , 
                 
                 8364
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010100; B = 7'b1110000; // Expected: {'P': 2240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010100; B = 7'b1110000; | Outputs: P=%b | Expected: P=%d",
                 1771,
                 
                 P
                 , 
                 
                 2240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011011; B = 7'b0111101; // Expected: {'P': 5551}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011011; B = 7'b0111101; | Outputs: P=%b | Expected: P=%d",
                 1772,
                 
                 P
                 , 
                 
                 5551
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111000; B = 7'b0011011; // Expected: {'P': 3240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111000; B = 7'b0011011; | Outputs: P=%b | Expected: P=%d",
                 1773,
                 
                 P
                 , 
                 
                 3240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100101; B = 7'b0100101; // Expected: {'P': 3737}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100101; B = 7'b0100101; | Outputs: P=%b | Expected: P=%d",
                 1774,
                 
                 P
                 , 
                 
                 3737
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110100; B = 7'b0000001; // Expected: {'P': 116}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110100; B = 7'b0000001; | Outputs: P=%b | Expected: P=%d",
                 1775,
                 
                 P
                 , 
                 
                 116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001000; B = 7'b1011111; // Expected: {'P': 6840}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001000; B = 7'b1011111; | Outputs: P=%b | Expected: P=%d",
                 1776,
                 
                 P
                 , 
                 
                 6840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010001; B = 7'b1001101; // Expected: {'P': 1309}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010001; B = 7'b1001101; | Outputs: P=%b | Expected: P=%d",
                 1777,
                 
                 P
                 , 
                 
                 1309
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111000; B = 7'b1110000; // Expected: {'P': 6272}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111000; B = 7'b1110000; | Outputs: P=%b | Expected: P=%d",
                 1778,
                 
                 P
                 , 
                 
                 6272
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101111; B = 7'b1001010; // Expected: {'P': 8214}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101111; B = 7'b1001010; | Outputs: P=%b | Expected: P=%d",
                 1779,
                 
                 P
                 , 
                 
                 8214
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001010; B = 7'b1110000; // Expected: {'P': 1120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001010; B = 7'b1110000; | Outputs: P=%b | Expected: P=%d",
                 1780,
                 
                 P
                 , 
                 
                 1120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011111; B = 7'b0111100; // Expected: {'P': 1860}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011111; B = 7'b0111100; | Outputs: P=%b | Expected: P=%d",
                 1781,
                 
                 P
                 , 
                 
                 1860
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110010; B = 7'b0111010; // Expected: {'P': 6612}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110010; B = 7'b0111010; | Outputs: P=%b | Expected: P=%d",
                 1782,
                 
                 P
                 , 
                 
                 6612
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001000; B = 7'b1000010; // Expected: {'P': 4752}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001000; B = 7'b1000010; | Outputs: P=%b | Expected: P=%d",
                 1783,
                 
                 P
                 , 
                 
                 4752
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010100; B = 7'b0000001; // Expected: {'P': 20}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010100; B = 7'b0000001; | Outputs: P=%b | Expected: P=%d",
                 1784,
                 
                 P
                 , 
                 
                 20
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110000; B = 7'b0100000; // Expected: {'P': 1536}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110000; B = 7'b0100000; | Outputs: P=%b | Expected: P=%d",
                 1785,
                 
                 P
                 , 
                 
                 1536
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101000; B = 7'b0000001; // Expected: {'P': 40}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101000; B = 7'b0000001; | Outputs: P=%b | Expected: P=%d",
                 1786,
                 
                 P
                 , 
                 
                 40
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100110; B = 7'b0001111; // Expected: {'P': 1530}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100110; B = 7'b0001111; | Outputs: P=%b | Expected: P=%d",
                 1787,
                 
                 P
                 , 
                 
                 1530
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111011; B = 7'b1010001; // Expected: {'P': 9963}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111011; B = 7'b1010001; | Outputs: P=%b | Expected: P=%d",
                 1788,
                 
                 P
                 , 
                 
                 9963
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001001; B = 7'b1000111; // Expected: {'P': 5183}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001001; B = 7'b1000111; | Outputs: P=%b | Expected: P=%d",
                 1789,
                 
                 P
                 , 
                 
                 5183
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011100; B = 7'b1011100; // Expected: {'P': 8464}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011100; B = 7'b1011100; | Outputs: P=%b | Expected: P=%d",
                 1790,
                 
                 P
                 , 
                 
                 8464
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010100; B = 7'b1101110; // Expected: {'P': 2200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010100; B = 7'b1101110; | Outputs: P=%b | Expected: P=%d",
                 1791,
                 
                 P
                 , 
                 
                 2200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100111; B = 7'b0100101; // Expected: {'P': 3811}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100111; B = 7'b0100101; | Outputs: P=%b | Expected: P=%d",
                 1792,
                 
                 P
                 , 
                 
                 3811
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011010; B = 7'b1001100; // Expected: {'P': 6840}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011010; B = 7'b1001100; | Outputs: P=%b | Expected: P=%d",
                 1793,
                 
                 P
                 , 
                 
                 6840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100001; B = 7'b0010000; // Expected: {'P': 528}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100001; B = 7'b0010000; | Outputs: P=%b | Expected: P=%d",
                 1794,
                 
                 P
                 , 
                 
                 528
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111011; B = 7'b1001111; // Expected: {'P': 4661}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111011; B = 7'b1001111; | Outputs: P=%b | Expected: P=%d",
                 1795,
                 
                 P
                 , 
                 
                 4661
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100111; B = 7'b1111000; // Expected: {'P': 4680}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100111; B = 7'b1111000; | Outputs: P=%b | Expected: P=%d",
                 1796,
                 
                 P
                 , 
                 
                 4680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001011; B = 7'b0110000; // Expected: {'P': 3600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001011; B = 7'b0110000; | Outputs: P=%b | Expected: P=%d",
                 1797,
                 
                 P
                 , 
                 
                 3600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000101; B = 7'b0001010; // Expected: {'P': 50}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000101; B = 7'b0001010; | Outputs: P=%b | Expected: P=%d",
                 1798,
                 
                 P
                 , 
                 
                 50
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101101; B = 7'b0000111; // Expected: {'P': 315}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101101; B = 7'b0000111; | Outputs: P=%b | Expected: P=%d",
                 1799,
                 
                 P
                 , 
                 
                 315
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010011; B = 7'b1111110; // Expected: {'P': 10458}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010011; B = 7'b1111110; | Outputs: P=%b | Expected: P=%d",
                 1800,
                 
                 P
                 , 
                 
                 10458
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110101; B = 7'b1011101; // Expected: {'P': 10881}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110101; B = 7'b1011101; | Outputs: P=%b | Expected: P=%d",
                 1801,
                 
                 P
                 , 
                 
                 10881
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000011; B = 7'b0100111; // Expected: {'P': 117}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000011; B = 7'b0100111; | Outputs: P=%b | Expected: P=%d",
                 1802,
                 
                 P
                 , 
                 
                 117
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101101; B = 7'b1101011; // Expected: {'P': 11663}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101101; B = 7'b1101011; | Outputs: P=%b | Expected: P=%d",
                 1803,
                 
                 P
                 , 
                 
                 11663
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001010; B = 7'b0011001; // Expected: {'P': 1850}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001010; B = 7'b0011001; | Outputs: P=%b | Expected: P=%d",
                 1804,
                 
                 P
                 , 
                 
                 1850
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101101; B = 7'b1001111; // Expected: {'P': 8611}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101101; B = 7'b1001111; | Outputs: P=%b | Expected: P=%d",
                 1805,
                 
                 P
                 , 
                 
                 8611
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001110; B = 7'b1100101; // Expected: {'P': 1414}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001110; B = 7'b1100101; | Outputs: P=%b | Expected: P=%d",
                 1806,
                 
                 P
                 , 
                 
                 1414
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011110; B = 7'b0111111; // Expected: {'P': 1890}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011110; B = 7'b0111111; | Outputs: P=%b | Expected: P=%d",
                 1807,
                 
                 P
                 , 
                 
                 1890
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100101; B = 7'b1100110; // Expected: {'P': 3774}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100101; B = 7'b1100110; | Outputs: P=%b | Expected: P=%d",
                 1808,
                 
                 P
                 , 
                 
                 3774
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101001; B = 7'b1101000; // Expected: {'P': 4264}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101001; B = 7'b1101000; | Outputs: P=%b | Expected: P=%d",
                 1809,
                 
                 P
                 , 
                 
                 4264
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111100; B = 7'b0100111; // Expected: {'P': 4836}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111100; B = 7'b0100111; | Outputs: P=%b | Expected: P=%d",
                 1810,
                 
                 P
                 , 
                 
                 4836
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010111; B = 7'b0110010; // Expected: {'P': 1150}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010111; B = 7'b0110010; | Outputs: P=%b | Expected: P=%d",
                 1811,
                 
                 P
                 , 
                 
                 1150
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101000; B = 7'b1011101; // Expected: {'P': 9672}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101000; B = 7'b1011101; | Outputs: P=%b | Expected: P=%d",
                 1812,
                 
                 P
                 , 
                 
                 9672
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000000; B = 7'b1000111; // Expected: {'P': 4544}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000000; B = 7'b1000111; | Outputs: P=%b | Expected: P=%d",
                 1813,
                 
                 P
                 , 
                 
                 4544
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001010; B = 7'b1110001; // Expected: {'P': 1130}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001010; B = 7'b1110001; | Outputs: P=%b | Expected: P=%d",
                 1814,
                 
                 P
                 , 
                 
                 1130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111110; B = 7'b1100001; // Expected: {'P': 12222}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111110; B = 7'b1100001; | Outputs: P=%b | Expected: P=%d",
                 1815,
                 
                 P
                 , 
                 
                 12222
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111100; B = 7'b0100010; // Expected: {'P': 2040}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111100; B = 7'b0100010; | Outputs: P=%b | Expected: P=%d",
                 1816,
                 
                 P
                 , 
                 
                 2040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011110; B = 7'b1010000; // Expected: {'P': 2400}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011110; B = 7'b1010000; | Outputs: P=%b | Expected: P=%d",
                 1817,
                 
                 P
                 , 
                 
                 2400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010000; B = 7'b1011100; // Expected: {'P': 7360}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010000; B = 7'b1011100; | Outputs: P=%b | Expected: P=%d",
                 1818,
                 
                 P
                 , 
                 
                 7360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011011; B = 7'b0101000; // Expected: {'P': 3640}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011011; B = 7'b0101000; | Outputs: P=%b | Expected: P=%d",
                 1819,
                 
                 P
                 , 
                 
                 3640
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001100; B = 7'b0011110; // Expected: {'P': 360}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001100; B = 7'b0011110; | Outputs: P=%b | Expected: P=%d",
                 1820,
                 
                 P
                 , 
                 
                 360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000111; B = 7'b0011010; // Expected: {'P': 182}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000111; B = 7'b0011010; | Outputs: P=%b | Expected: P=%d",
                 1821,
                 
                 P
                 , 
                 
                 182
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100101; B = 7'b1010001; // Expected: {'P': 8181}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100101; B = 7'b1010001; | Outputs: P=%b | Expected: P=%d",
                 1822,
                 
                 P
                 , 
                 
                 8181
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010000; B = 7'b1011010; // Expected: {'P': 7200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010000; B = 7'b1011010; | Outputs: P=%b | Expected: P=%d",
                 1823,
                 
                 P
                 , 
                 
                 7200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110110; B = 7'b1100010; // Expected: {'P': 5292}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110110; B = 7'b1100010; | Outputs: P=%b | Expected: P=%d",
                 1824,
                 
                 P
                 , 
                 
                 5292
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001000; B = 7'b0000100; // Expected: {'P': 288}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001000; B = 7'b0000100; | Outputs: P=%b | Expected: P=%d",
                 1825,
                 
                 P
                 , 
                 
                 288
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011111; B = 7'b1101010; // Expected: {'P': 3286}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011111; B = 7'b1101010; | Outputs: P=%b | Expected: P=%d",
                 1826,
                 
                 P
                 , 
                 
                 3286
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101111; B = 7'b0100101; // Expected: {'P': 4107}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101111; B = 7'b0100101; | Outputs: P=%b | Expected: P=%d",
                 1827,
                 
                 P
                 , 
                 
                 4107
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001000; B = 7'b1001110; // Expected: {'P': 5616}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001000; B = 7'b1001110; | Outputs: P=%b | Expected: P=%d",
                 1828,
                 
                 P
                 , 
                 
                 5616
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111111; B = 7'b0100111; // Expected: {'P': 4953}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111111; B = 7'b0100111; | Outputs: P=%b | Expected: P=%d",
                 1829,
                 
                 P
                 , 
                 
                 4953
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101111; B = 7'b1001101; // Expected: {'P': 8547}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101111; B = 7'b1001101; | Outputs: P=%b | Expected: P=%d",
                 1830,
                 
                 P
                 , 
                 
                 8547
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101100; B = 7'b0011110; // Expected: {'P': 3240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101100; B = 7'b0011110; | Outputs: P=%b | Expected: P=%d",
                 1831,
                 
                 P
                 , 
                 
                 3240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010001; B = 7'b0011001; // Expected: {'P': 2025}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010001; B = 7'b0011001; | Outputs: P=%b | Expected: P=%d",
                 1832,
                 
                 P
                 , 
                 
                 2025
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000111; B = 7'b0111110; // Expected: {'P': 434}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000111; B = 7'b0111110; | Outputs: P=%b | Expected: P=%d",
                 1833,
                 
                 P
                 , 
                 
                 434
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110001; B = 7'b0110110; // Expected: {'P': 2646}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110001; B = 7'b0110110; | Outputs: P=%b | Expected: P=%d",
                 1834,
                 
                 P
                 , 
                 
                 2646
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110010; B = 7'b1110110; // Expected: {'P': 5900}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110010; B = 7'b1110110; | Outputs: P=%b | Expected: P=%d",
                 1835,
                 
                 P
                 , 
                 
                 5900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011101; B = 7'b1111001; // Expected: {'P': 3509}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011101; B = 7'b1111001; | Outputs: P=%b | Expected: P=%d",
                 1836,
                 
                 P
                 , 
                 
                 3509
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101111; B = 7'b0101000; // Expected: {'P': 4440}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101111; B = 7'b0101000; | Outputs: P=%b | Expected: P=%d",
                 1837,
                 
                 P
                 , 
                 
                 4440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101111; B = 7'b0010001; // Expected: {'P': 799}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101111; B = 7'b0010001; | Outputs: P=%b | Expected: P=%d",
                 1838,
                 
                 P
                 , 
                 
                 799
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000110; B = 7'b0011000; // Expected: {'P': 1680}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000110; B = 7'b0011000; | Outputs: P=%b | Expected: P=%d",
                 1839,
                 
                 P
                 , 
                 
                 1680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110010; B = 7'b1011100; // Expected: {'P': 10488}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110010; B = 7'b1011100; | Outputs: P=%b | Expected: P=%d",
                 1840,
                 
                 P
                 , 
                 
                 10488
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111110; B = 7'b1001011; // Expected: {'P': 9450}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111110; B = 7'b1001011; | Outputs: P=%b | Expected: P=%d",
                 1841,
                 
                 P
                 , 
                 
                 9450
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001001; B = 7'b0000101; // Expected: {'P': 365}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001001; B = 7'b0000101; | Outputs: P=%b | Expected: P=%d",
                 1842,
                 
                 P
                 , 
                 
                 365
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001111; B = 7'b0101000; // Expected: {'P': 600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001111; B = 7'b0101000; | Outputs: P=%b | Expected: P=%d",
                 1843,
                 
                 P
                 , 
                 
                 600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110110; B = 7'b1101000; // Expected: {'P': 5616}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110110; B = 7'b1101000; | Outputs: P=%b | Expected: P=%d",
                 1844,
                 
                 P
                 , 
                 
                 5616
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011101; B = 7'b0100101; // Expected: {'P': 1073}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011101; B = 7'b0100101; | Outputs: P=%b | Expected: P=%d",
                 1845,
                 
                 P
                 , 
                 
                 1073
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010001; B = 7'b1011000; // Expected: {'P': 1496}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010001; B = 7'b1011000; | Outputs: P=%b | Expected: P=%d",
                 1846,
                 
                 P
                 , 
                 
                 1496
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001001; B = 7'b0101100; // Expected: {'P': 396}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001001; B = 7'b0101100; | Outputs: P=%b | Expected: P=%d",
                 1847,
                 
                 P
                 , 
                 
                 396
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001100; B = 7'b1110100; // Expected: {'P': 8816}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001100; B = 7'b1110100; | Outputs: P=%b | Expected: P=%d",
                 1848,
                 
                 P
                 , 
                 
                 8816
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010000; B = 7'b1011011; // Expected: {'P': 1456}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010000; B = 7'b1011011; | Outputs: P=%b | Expected: P=%d",
                 1849,
                 
                 P
                 , 
                 
                 1456
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000000; B = 7'b1110100; // Expected: {'P': 7424}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000000; B = 7'b1110100; | Outputs: P=%b | Expected: P=%d",
                 1850,
                 
                 P
                 , 
                 
                 7424
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001010; B = 7'b1001100; // Expected: {'P': 760}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001010; B = 7'b1001100; | Outputs: P=%b | Expected: P=%d",
                 1851,
                 
                 P
                 , 
                 
                 760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000011; B = 7'b0010110; // Expected: {'P': 1474}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000011; B = 7'b0010110; | Outputs: P=%b | Expected: P=%d",
                 1852,
                 
                 P
                 , 
                 
                 1474
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001011; B = 7'b1000111; // Expected: {'P': 781}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001011; B = 7'b1000111; | Outputs: P=%b | Expected: P=%d",
                 1853,
                 
                 P
                 , 
                 
                 781
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001000; B = 7'b1001100; // Expected: {'P': 5472}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001000; B = 7'b1001100; | Outputs: P=%b | Expected: P=%d",
                 1854,
                 
                 P
                 , 
                 
                 5472
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001110; B = 7'b1000010; // Expected: {'P': 5148}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001110; B = 7'b1000010; | Outputs: P=%b | Expected: P=%d",
                 1855,
                 
                 P
                 , 
                 
                 5148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100100; B = 7'b0010110; // Expected: {'P': 792}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100100; B = 7'b0010110; | Outputs: P=%b | Expected: P=%d",
                 1856,
                 
                 P
                 , 
                 
                 792
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001110; B = 7'b1011010; // Expected: {'P': 7020}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001110; B = 7'b1011010; | Outputs: P=%b | Expected: P=%d",
                 1857,
                 
                 P
                 , 
                 
                 7020
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110001; B = 7'b0100100; // Expected: {'P': 4068}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110001; B = 7'b0100100; | Outputs: P=%b | Expected: P=%d",
                 1858,
                 
                 P
                 , 
                 
                 4068
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101001; B = 7'b0001010; // Expected: {'P': 410}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101001; B = 7'b0001010; | Outputs: P=%b | Expected: P=%d",
                 1859,
                 
                 P
                 , 
                 
                 410
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011101; B = 7'b1111001; // Expected: {'P': 11253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011101; B = 7'b1111001; | Outputs: P=%b | Expected: P=%d",
                 1860,
                 
                 P
                 , 
                 
                 11253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010101; B = 7'b1011011; // Expected: {'P': 1911}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010101; B = 7'b1011011; | Outputs: P=%b | Expected: P=%d",
                 1861,
                 
                 P
                 , 
                 
                 1911
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101000; B = 7'b0100011; // Expected: {'P': 1400}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101000; B = 7'b0100011; | Outputs: P=%b | Expected: P=%d",
                 1862,
                 
                 P
                 , 
                 
                 1400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111110; B = 7'b1111000; // Expected: {'P': 7440}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111110; B = 7'b1111000; | Outputs: P=%b | Expected: P=%d",
                 1863,
                 
                 P
                 , 
                 
                 7440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011111; B = 7'b1000010; // Expected: {'P': 6270}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011111; B = 7'b1000010; | Outputs: P=%b | Expected: P=%d",
                 1864,
                 
                 P
                 , 
                 
                 6270
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000011; B = 7'b0100011; // Expected: {'P': 2345}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000011; B = 7'b0100011; | Outputs: P=%b | Expected: P=%d",
                 1865,
                 
                 P
                 , 
                 
                 2345
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011111; B = 7'b1111100; // Expected: {'P': 11780}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011111; B = 7'b1111100; | Outputs: P=%b | Expected: P=%d",
                 1866,
                 
                 P
                 , 
                 
                 11780
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101011; B = 7'b1100100; // Expected: {'P': 10700}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101011; B = 7'b1100100; | Outputs: P=%b | Expected: P=%d",
                 1867,
                 
                 P
                 , 
                 
                 10700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111011; B = 7'b1111011; // Expected: {'P': 7257}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111011; B = 7'b1111011; | Outputs: P=%b | Expected: P=%d",
                 1868,
                 
                 P
                 , 
                 
                 7257
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010011; B = 7'b0010100; // Expected: {'P': 1660}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010011; B = 7'b0010100; | Outputs: P=%b | Expected: P=%d",
                 1869,
                 
                 P
                 , 
                 
                 1660
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101001; B = 7'b0011010; // Expected: {'P': 1066}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101001; B = 7'b0011010; | Outputs: P=%b | Expected: P=%d",
                 1870,
                 
                 P
                 , 
                 
                 1066
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001110; B = 7'b1011001; // Expected: {'P': 1246}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001110; B = 7'b1011001; | Outputs: P=%b | Expected: P=%d",
                 1871,
                 
                 P
                 , 
                 
                 1246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101001; B = 7'b1011001; // Expected: {'P': 3649}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101001; B = 7'b1011001; | Outputs: P=%b | Expected: P=%d",
                 1872,
                 
                 P
                 , 
                 
                 3649
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001111; B = 7'b1101110; // Expected: {'P': 8690}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001111; B = 7'b1101110; | Outputs: P=%b | Expected: P=%d",
                 1873,
                 
                 P
                 , 
                 
                 8690
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011000; B = 7'b0010100; // Expected: {'P': 480}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011000; B = 7'b0010100; | Outputs: P=%b | Expected: P=%d",
                 1874,
                 
                 P
                 , 
                 
                 480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111100; B = 7'b0111111; // Expected: {'P': 7812}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111100; B = 7'b0111111; | Outputs: P=%b | Expected: P=%d",
                 1875,
                 
                 P
                 , 
                 
                 7812
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110000; B = 7'b0001001; // Expected: {'P': 1008}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110000; B = 7'b0001001; | Outputs: P=%b | Expected: P=%d",
                 1876,
                 
                 P
                 , 
                 
                 1008
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001100; B = 7'b1000100; // Expected: {'P': 5168}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001100; B = 7'b1000100; | Outputs: P=%b | Expected: P=%d",
                 1877,
                 
                 P
                 , 
                 
                 5168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011111; B = 7'b0100101; // Expected: {'P': 3515}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011111; B = 7'b0100101; | Outputs: P=%b | Expected: P=%d",
                 1878,
                 
                 P
                 , 
                 
                 3515
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110010; B = 7'b0010100; // Expected: {'P': 2280}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110010; B = 7'b0010100; | Outputs: P=%b | Expected: P=%d",
                 1879,
                 
                 P
                 , 
                 
                 2280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110111; B = 7'b1001101; // Expected: {'P': 9163}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110111; B = 7'b1001101; | Outputs: P=%b | Expected: P=%d",
                 1880,
                 
                 P
                 , 
                 
                 9163
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100010; B = 7'b0000111; // Expected: {'P': 238}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100010; B = 7'b0000111; | Outputs: P=%b | Expected: P=%d",
                 1881,
                 
                 P
                 , 
                 
                 238
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110101; B = 7'b0010101; // Expected: {'P': 1113}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110101; B = 7'b0010101; | Outputs: P=%b | Expected: P=%d",
                 1882,
                 
                 P
                 , 
                 
                 1113
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111010; B = 7'b1000000; // Expected: {'P': 7808}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111010; B = 7'b1000000; | Outputs: P=%b | Expected: P=%d",
                 1883,
                 
                 P
                 , 
                 
                 7808
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001110; B = 7'b1000000; // Expected: {'P': 896}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001110; B = 7'b1000000; | Outputs: P=%b | Expected: P=%d",
                 1884,
                 
                 P
                 , 
                 
                 896
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000010; B = 7'b0111100; // Expected: {'P': 3960}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000010; B = 7'b0111100; | Outputs: P=%b | Expected: P=%d",
                 1885,
                 
                 P
                 , 
                 
                 3960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010000; B = 7'b0011110; // Expected: {'P': 2400}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010000; B = 7'b0011110; | Outputs: P=%b | Expected: P=%d",
                 1886,
                 
                 P
                 , 
                 
                 2400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111010; B = 7'b1111110; // Expected: {'P': 15372}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111010; B = 7'b1111110; | Outputs: P=%b | Expected: P=%d",
                 1887,
                 
                 P
                 , 
                 
                 15372
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011010; B = 7'b0111110; // Expected: {'P': 5580}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011010; B = 7'b0111110; | Outputs: P=%b | Expected: P=%d",
                 1888,
                 
                 P
                 , 
                 
                 5580
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010100; B = 7'b1000011; // Expected: {'P': 5628}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010100; B = 7'b1000011; | Outputs: P=%b | Expected: P=%d",
                 1889,
                 
                 P
                 , 
                 
                 5628
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111111; B = 7'b0110111; // Expected: {'P': 6985}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111111; B = 7'b0110111; | Outputs: P=%b | Expected: P=%d",
                 1890,
                 
                 P
                 , 
                 
                 6985
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100100; B = 7'b1000001; // Expected: {'P': 6500}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100100; B = 7'b1000001; | Outputs: P=%b | Expected: P=%d",
                 1891,
                 
                 P
                 , 
                 
                 6500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111001; B = 7'b0100111; // Expected: {'P': 2223}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111001; B = 7'b0100111; | Outputs: P=%b | Expected: P=%d",
                 1892,
                 
                 P
                 , 
                 
                 2223
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101101; B = 7'b0100011; // Expected: {'P': 3815}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101101; B = 7'b0100011; | Outputs: P=%b | Expected: P=%d",
                 1893,
                 
                 P
                 , 
                 
                 3815
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011111; B = 7'b1001010; // Expected: {'P': 7030}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011111; B = 7'b1001010; | Outputs: P=%b | Expected: P=%d",
                 1894,
                 
                 P
                 , 
                 
                 7030
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000100; B = 7'b0100011; // Expected: {'P': 140}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000100; B = 7'b0100011; | Outputs: P=%b | Expected: P=%d",
                 1895,
                 
                 P
                 , 
                 
                 140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111001; B = 7'b0111100; // Expected: {'P': 7260}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111001; B = 7'b0111100; | Outputs: P=%b | Expected: P=%d",
                 1896,
                 
                 P
                 , 
                 
                 7260
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001111; B = 7'b0011110; // Expected: {'P': 2370}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001111; B = 7'b0011110; | Outputs: P=%b | Expected: P=%d",
                 1897,
                 
                 P
                 , 
                 
                 2370
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001001; B = 7'b0010010; // Expected: {'P': 162}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001001; B = 7'b0010010; | Outputs: P=%b | Expected: P=%d",
                 1898,
                 
                 P
                 , 
                 
                 162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110000; B = 7'b1000000; // Expected: {'P': 7168}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110000; B = 7'b1000000; | Outputs: P=%b | Expected: P=%d",
                 1899,
                 
                 P
                 , 
                 
                 7168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111111; B = 7'b0110110; // Expected: {'P': 3402}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111111; B = 7'b0110110; | Outputs: P=%b | Expected: P=%d",
                 1900,
                 
                 P
                 , 
                 
                 3402
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010110; B = 7'b1001011; // Expected: {'P': 1650}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010110; B = 7'b1001011; | Outputs: P=%b | Expected: P=%d",
                 1901,
                 
                 P
                 , 
                 
                 1650
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110101; B = 7'b0111111; // Expected: {'P': 3339}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110101; B = 7'b0111111; | Outputs: P=%b | Expected: P=%d",
                 1902,
                 
                 P
                 , 
                 
                 3339
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000101; B = 7'b0010100; // Expected: {'P': 1380}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000101; B = 7'b0010100; | Outputs: P=%b | Expected: P=%d",
                 1903,
                 
                 P
                 , 
                 
                 1380
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010111; B = 7'b1001110; // Expected: {'P': 1794}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010111; B = 7'b1001110; | Outputs: P=%b | Expected: P=%d",
                 1904,
                 
                 P
                 , 
                 
                 1794
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010111; B = 7'b1001001; // Expected: {'P': 6351}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010111; B = 7'b1001001; | Outputs: P=%b | Expected: P=%d",
                 1905,
                 
                 P
                 , 
                 
                 6351
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110111; B = 7'b1000001; // Expected: {'P': 3575}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110111; B = 7'b1000001; | Outputs: P=%b | Expected: P=%d",
                 1906,
                 
                 P
                 , 
                 
                 3575
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011001; B = 7'b0001010; // Expected: {'P': 890}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011001; B = 7'b0001010; | Outputs: P=%b | Expected: P=%d",
                 1907,
                 
                 P
                 , 
                 
                 890
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100110; B = 7'b0000001; // Expected: {'P': 38}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100110; B = 7'b0000001; | Outputs: P=%b | Expected: P=%d",
                 1908,
                 
                 P
                 , 
                 
                 38
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011100; B = 7'b0001100; // Expected: {'P': 1104}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011100; B = 7'b0001100; | Outputs: P=%b | Expected: P=%d",
                 1909,
                 
                 P
                 , 
                 
                 1104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100011; B = 7'b1000100; // Expected: {'P': 2380}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100011; B = 7'b1000100; | Outputs: P=%b | Expected: P=%d",
                 1910,
                 
                 P
                 , 
                 
                 2380
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100111; B = 7'b0110111; // Expected: {'P': 2145}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100111; B = 7'b0110111; | Outputs: P=%b | Expected: P=%d",
                 1911,
                 
                 P
                 , 
                 
                 2145
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101001; B = 7'b0001100; // Expected: {'P': 492}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101001; B = 7'b0001100; | Outputs: P=%b | Expected: P=%d",
                 1912,
                 
                 P
                 , 
                 
                 492
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011011; B = 7'b0101100; // Expected: {'P': 4004}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011011; B = 7'b0101100; | Outputs: P=%b | Expected: P=%d",
                 1913,
                 
                 P
                 , 
                 
                 4004
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001110; B = 7'b0010100; // Expected: {'P': 280}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001110; B = 7'b0010100; | Outputs: P=%b | Expected: P=%d",
                 1914,
                 
                 P
                 , 
                 
                 280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101100; B = 7'b0000100; // Expected: {'P': 176}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101100; B = 7'b0000100; | Outputs: P=%b | Expected: P=%d",
                 1915,
                 
                 P
                 , 
                 
                 176
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101111; B = 7'b1110010; // Expected: {'P': 12654}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101111; B = 7'b1110010; | Outputs: P=%b | Expected: P=%d",
                 1916,
                 
                 P
                 , 
                 
                 12654
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000100; B = 7'b0011110; // Expected: {'P': 2040}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000100; B = 7'b0011110; | Outputs: P=%b | Expected: P=%d",
                 1917,
                 
                 P
                 , 
                 
                 2040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111011; B = 7'b1110000; // Expected: {'P': 13776}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111011; B = 7'b1110000; | Outputs: P=%b | Expected: P=%d",
                 1918,
                 
                 P
                 , 
                 
                 13776
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111101; B = 7'b0001100; // Expected: {'P': 732}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111101; B = 7'b0001100; | Outputs: P=%b | Expected: P=%d",
                 1919,
                 
                 P
                 , 
                 
                 732
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101001; B = 7'b0111111; // Expected: {'P': 6615}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101001; B = 7'b0111111; | Outputs: P=%b | Expected: P=%d",
                 1920,
                 
                 P
                 , 
                 
                 6615
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011010; B = 7'b0010001; // Expected: {'P': 442}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011010; B = 7'b0010001; | Outputs: P=%b | Expected: P=%d",
                 1921,
                 
                 P
                 , 
                 
                 442
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100000; B = 7'b0000100; // Expected: {'P': 128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100000; B = 7'b0000100; | Outputs: P=%b | Expected: P=%d",
                 1922,
                 
                 P
                 , 
                 
                 128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110011; B = 7'b1100111; // Expected: {'P': 5253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110011; B = 7'b1100111; | Outputs: P=%b | Expected: P=%d",
                 1923,
                 
                 P
                 , 
                 
                 5253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001111; B = 7'b1001010; // Expected: {'P': 1110}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001111; B = 7'b1001010; | Outputs: P=%b | Expected: P=%d",
                 1924,
                 
                 P
                 , 
                 
                 1110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010110; B = 7'b1010101; // Expected: {'P': 1870}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010110; B = 7'b1010101; | Outputs: P=%b | Expected: P=%d",
                 1925,
                 
                 P
                 , 
                 
                 1870
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000111; B = 7'b0100110; // Expected: {'P': 266}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000111; B = 7'b0100110; | Outputs: P=%b | Expected: P=%d",
                 1926,
                 
                 P
                 , 
                 
                 266
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101101; B = 7'b1110011; // Expected: {'P': 5175}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101101; B = 7'b1110011; | Outputs: P=%b | Expected: P=%d",
                 1927,
                 
                 P
                 , 
                 
                 5175
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010001; B = 7'b1000000; // Expected: {'P': 1088}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010001; B = 7'b1000000; | Outputs: P=%b | Expected: P=%d",
                 1928,
                 
                 P
                 , 
                 
                 1088
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110000; B = 7'b0111110; // Expected: {'P': 6944}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110000; B = 7'b0111110; | Outputs: P=%b | Expected: P=%d",
                 1929,
                 
                 P
                 , 
                 
                 6944
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111010; B = 7'b1001100; // Expected: {'P': 9272}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111010; B = 7'b1001100; | Outputs: P=%b | Expected: P=%d",
                 1930,
                 
                 P
                 , 
                 
                 9272
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100111; B = 7'b1100011; // Expected: {'P': 10197}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100111; B = 7'b1100011; | Outputs: P=%b | Expected: P=%d",
                 1931,
                 
                 P
                 , 
                 
                 10197
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011010; B = 7'b1100001; // Expected: {'P': 2522}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011010; B = 7'b1100001; | Outputs: P=%b | Expected: P=%d",
                 1932,
                 
                 P
                 , 
                 
                 2522
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101001; B = 7'b1100100; // Expected: {'P': 4100}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101001; B = 7'b1100100; | Outputs: P=%b | Expected: P=%d",
                 1933,
                 
                 P
                 , 
                 
                 4100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101010; B = 7'b0100010; // Expected: {'P': 3604}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101010; B = 7'b0100010; | Outputs: P=%b | Expected: P=%d",
                 1934,
                 
                 P
                 , 
                 
                 3604
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001111; B = 7'b1011011; // Expected: {'P': 7189}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001111; B = 7'b1011011; | Outputs: P=%b | Expected: P=%d",
                 1935,
                 
                 P
                 , 
                 
                 7189
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100111; B = 7'b0001000; // Expected: {'P': 824}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100111; B = 7'b0001000; | Outputs: P=%b | Expected: P=%d",
                 1936,
                 
                 P
                 , 
                 
                 824
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101010; B = 7'b0010001; // Expected: {'P': 714}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101010; B = 7'b0010001; | Outputs: P=%b | Expected: P=%d",
                 1937,
                 
                 P
                 , 
                 
                 714
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010111; B = 7'b1010000; // Expected: {'P': 6960}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010111; B = 7'b1010000; | Outputs: P=%b | Expected: P=%d",
                 1938,
                 
                 P
                 , 
                 
                 6960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111110; B = 7'b1011100; // Expected: {'P': 5704}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111110; B = 7'b1011100; | Outputs: P=%b | Expected: P=%d",
                 1939,
                 
                 P
                 , 
                 
                 5704
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010100; B = 7'b0101000; // Expected: {'P': 800}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010100; B = 7'b0101000; | Outputs: P=%b | Expected: P=%d",
                 1940,
                 
                 P
                 , 
                 
                 800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110010; B = 7'b1011111; // Expected: {'P': 10830}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110010; B = 7'b1011111; | Outputs: P=%b | Expected: P=%d",
                 1941,
                 
                 P
                 , 
                 
                 10830
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001111; B = 7'b0110101; // Expected: {'P': 795}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001111; B = 7'b0110101; | Outputs: P=%b | Expected: P=%d",
                 1942,
                 
                 P
                 , 
                 
                 795
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100011; B = 7'b0110101; // Expected: {'P': 5247}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100011; B = 7'b0110101; | Outputs: P=%b | Expected: P=%d",
                 1943,
                 
                 P
                 , 
                 
                 5247
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110001; B = 7'b0100101; // Expected: {'P': 1813}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110001; B = 7'b0100101; | Outputs: P=%b | Expected: P=%d",
                 1944,
                 
                 P
                 , 
                 
                 1813
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010100; B = 7'b0101011; // Expected: {'P': 860}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010100; B = 7'b0101011; | Outputs: P=%b | Expected: P=%d",
                 1945,
                 
                 P
                 , 
                 
                 860
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000100; B = 7'b0100111; // Expected: {'P': 156}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000100; B = 7'b0100111; | Outputs: P=%b | Expected: P=%d",
                 1946,
                 
                 P
                 , 
                 
                 156
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001111; B = 7'b0111100; // Expected: {'P': 900}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001111; B = 7'b0111100; | Outputs: P=%b | Expected: P=%d",
                 1947,
                 
                 P
                 , 
                 
                 900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101000; B = 7'b0001011; // Expected: {'P': 440}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101000; B = 7'b0001011; | Outputs: P=%b | Expected: P=%d",
                 1948,
                 
                 P
                 , 
                 
                 440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101001; B = 7'b1001110; // Expected: {'P': 8190}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101001; B = 7'b1001110; | Outputs: P=%b | Expected: P=%d",
                 1949,
                 
                 P
                 , 
                 
                 8190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001110; B = 7'b0110101; // Expected: {'P': 742}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001110; B = 7'b0110101; | Outputs: P=%b | Expected: P=%d",
                 1950,
                 
                 P
                 , 
                 
                 742
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110110; B = 7'b1111000; // Expected: {'P': 6480}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110110; B = 7'b1111000; | Outputs: P=%b | Expected: P=%d",
                 1951,
                 
                 P
                 , 
                 
                 6480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110101; B = 7'b0110000; // Expected: {'P': 2544}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110101; B = 7'b0110000; | Outputs: P=%b | Expected: P=%d",
                 1952,
                 
                 P
                 , 
                 
                 2544
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101100; B = 7'b1101001; // Expected: {'P': 4620}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101100; B = 7'b1101001; | Outputs: P=%b | Expected: P=%d",
                 1953,
                 
                 P
                 , 
                 
                 4620
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110101; B = 7'b0001010; // Expected: {'P': 530}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110101; B = 7'b0001010; | Outputs: P=%b | Expected: P=%d",
                 1954,
                 
                 P
                 , 
                 
                 530
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000110; B = 7'b1110000; // Expected: {'P': 672}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000110; B = 7'b1110000; | Outputs: P=%b | Expected: P=%d",
                 1955,
                 
                 P
                 , 
                 
                 672
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011001; B = 7'b0101101; // Expected: {'P': 1125}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011001; B = 7'b0101101; | Outputs: P=%b | Expected: P=%d",
                 1956,
                 
                 P
                 , 
                 
                 1125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000010; B = 7'b1101111; // Expected: {'P': 222}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000010; B = 7'b1101111; | Outputs: P=%b | Expected: P=%d",
                 1957,
                 
                 P
                 , 
                 
                 222
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011000; B = 7'b1001100; // Expected: {'P': 6688}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011000; B = 7'b1001100; | Outputs: P=%b | Expected: P=%d",
                 1958,
                 
                 P
                 , 
                 
                 6688
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101111; B = 7'b1001111; // Expected: {'P': 8769}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101111; B = 7'b1001111; | Outputs: P=%b | Expected: P=%d",
                 1959,
                 
                 P
                 , 
                 
                 8769
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110111; B = 7'b0001000; // Expected: {'P': 952}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110111; B = 7'b0001000; | Outputs: P=%b | Expected: P=%d",
                 1960,
                 
                 P
                 , 
                 
                 952
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011110; B = 7'b1101110; // Expected: {'P': 10340}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011110; B = 7'b1101110; | Outputs: P=%b | Expected: P=%d",
                 1961,
                 
                 P
                 , 
                 
                 10340
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010001; B = 7'b1000001; // Expected: {'P': 5265}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010001; B = 7'b1000001; | Outputs: P=%b | Expected: P=%d",
                 1962,
                 
                 P
                 , 
                 
                 5265
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100000; B = 7'b1000110; // Expected: {'P': 2240}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100000; B = 7'b1000110; | Outputs: P=%b | Expected: P=%d",
                 1963,
                 
                 P
                 , 
                 
                 2240
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001101; B = 7'b0010111; // Expected: {'P': 1771}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001101; B = 7'b0010111; | Outputs: P=%b | Expected: P=%d",
                 1964,
                 
                 P
                 , 
                 
                 1771
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001100; B = 7'b1011011; // Expected: {'P': 1092}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001100; B = 7'b1011011; | Outputs: P=%b | Expected: P=%d",
                 1965,
                 
                 P
                 , 
                 
                 1092
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100111; B = 7'b0000100; // Expected: {'P': 412}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100111; B = 7'b0000100; | Outputs: P=%b | Expected: P=%d",
                 1966,
                 
                 P
                 , 
                 
                 412
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101011; B = 7'b1011101; // Expected: {'P': 9951}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101011; B = 7'b1011101; | Outputs: P=%b | Expected: P=%d",
                 1967,
                 
                 P
                 , 
                 
                 9951
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010111; B = 7'b0000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010111; B = 7'b0000000; | Outputs: P=%b | Expected: P=%d",
                 1968,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100100; B = 7'b1101001; // Expected: {'P': 3780}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100100; B = 7'b1101001; | Outputs: P=%b | Expected: P=%d",
                 1969,
                 
                 P
                 , 
                 
                 3780
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000111; B = 7'b1011100; // Expected: {'P': 6532}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000111; B = 7'b1011100; | Outputs: P=%b | Expected: P=%d",
                 1970,
                 
                 P
                 , 
                 
                 6532
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000000; B = 7'b1010010; // Expected: {'P': 5248}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000000; B = 7'b1010010; | Outputs: P=%b | Expected: P=%d",
                 1971,
                 
                 P
                 , 
                 
                 5248
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101101; B = 7'b0110101; // Expected: {'P': 2385}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101101; B = 7'b0110101; | Outputs: P=%b | Expected: P=%d",
                 1972,
                 
                 P
                 , 
                 
                 2385
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110011; B = 7'b0011101; // Expected: {'P': 1479}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110011; B = 7'b0011101; | Outputs: P=%b | Expected: P=%d",
                 1973,
                 
                 P
                 , 
                 
                 1479
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100100; B = 7'b0111111; // Expected: {'P': 6300}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100100; B = 7'b0111111; | Outputs: P=%b | Expected: P=%d",
                 1974,
                 
                 P
                 , 
                 
                 6300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001101; B = 7'b1101101; // Expected: {'P': 1417}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001101; B = 7'b1101101; | Outputs: P=%b | Expected: P=%d",
                 1975,
                 
                 P
                 , 
                 
                 1417
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101010; B = 7'b1111010; // Expected: {'P': 12932}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101010; B = 7'b1111010; | Outputs: P=%b | Expected: P=%d",
                 1976,
                 
                 P
                 , 
                 
                 12932
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111010; B = 7'b0111011; // Expected: {'P': 7198}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111010; B = 7'b0111011; | Outputs: P=%b | Expected: P=%d",
                 1977,
                 
                 P
                 , 
                 
                 7198
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111011; B = 7'b0111110; // Expected: {'P': 3658}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111011; B = 7'b0111110; | Outputs: P=%b | Expected: P=%d",
                 1978,
                 
                 P
                 , 
                 
                 3658
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000100; B = 7'b0011001; // Expected: {'P': 1700}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000100; B = 7'b0011001; | Outputs: P=%b | Expected: P=%d",
                 1979,
                 
                 P
                 , 
                 
                 1700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000000; B = 7'b1110010; // Expected: {'P': 7296}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000000; B = 7'b1110010; | Outputs: P=%b | Expected: P=%d",
                 1980,
                 
                 P
                 , 
                 
                 7296
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010010; B = 7'b0010010; // Expected: {'P': 324}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010010; B = 7'b0010010; | Outputs: P=%b | Expected: P=%d",
                 1981,
                 
                 P
                 , 
                 
                 324
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111110; B = 7'b0101111; // Expected: {'P': 5922}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111110; B = 7'b0101111; | Outputs: P=%b | Expected: P=%d",
                 1982,
                 
                 P
                 , 
                 
                 5922
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010111; B = 7'b0110110; // Expected: {'P': 4698}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010111; B = 7'b0110110; | Outputs: P=%b | Expected: P=%d",
                 1983,
                 
                 P
                 , 
                 
                 4698
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101110; B = 7'b1011100; // Expected: {'P': 10120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101110; B = 7'b1011100; | Outputs: P=%b | Expected: P=%d",
                 1984,
                 
                 P
                 , 
                 
                 10120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000000; B = 7'b0011001; // Expected: {'P': 1600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000000; B = 7'b0011001; | Outputs: P=%b | Expected: P=%d",
                 1985,
                 
                 P
                 , 
                 
                 1600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100111; B = 7'b0000110; // Expected: {'P': 234}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100111; B = 7'b0000110; | Outputs: P=%b | Expected: P=%d",
                 1986,
                 
                 P
                 , 
                 
                 234
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011011; B = 7'b0001000; // Expected: {'P': 216}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011011; B = 7'b0001000; | Outputs: P=%b | Expected: P=%d",
                 1987,
                 
                 P
                 , 
                 
                 216
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111000; B = 7'b1000000; // Expected: {'P': 7680}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111000; B = 7'b1000000; | Outputs: P=%b | Expected: P=%d",
                 1988,
                 
                 P
                 , 
                 
                 7680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010011; B = 7'b0111110; // Expected: {'P': 1178}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010011; B = 7'b0111110; | Outputs: P=%b | Expected: P=%d",
                 1989,
                 
                 P
                 , 
                 
                 1178
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010010; B = 7'b1111101; // Expected: {'P': 2250}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010010; B = 7'b1111101; | Outputs: P=%b | Expected: P=%d",
                 1990,
                 
                 P
                 , 
                 
                 2250
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100111; B = 7'b0001100; // Expected: {'P': 1236}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100111; B = 7'b0001100; | Outputs: P=%b | Expected: P=%d",
                 1991,
                 
                 P
                 , 
                 
                 1236
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001010; B = 7'b1101111; // Expected: {'P': 1110}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001010; B = 7'b1101111; | Outputs: P=%b | Expected: P=%d",
                 1992,
                 
                 P
                 , 
                 
                 1110
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101100; B = 7'b0111101; // Expected: {'P': 6588}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101100; B = 7'b0111101; | Outputs: P=%b | Expected: P=%d",
                 1993,
                 
                 P
                 , 
                 
                 6588
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110110; B = 7'b0101001; // Expected: {'P': 2214}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110110; B = 7'b0101001; | Outputs: P=%b | Expected: P=%d",
                 1994,
                 
                 P
                 , 
                 
                 2214
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001010; B = 7'b0100111; // Expected: {'P': 2886}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001010; B = 7'b0100111; | Outputs: P=%b | Expected: P=%d",
                 1995,
                 
                 P
                 , 
                 
                 2886
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111110; B = 7'b0110111; // Expected: {'P': 3410}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111110; B = 7'b0110111; | Outputs: P=%b | Expected: P=%d",
                 1996,
                 
                 P
                 , 
                 
                 3410
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100001; B = 7'b0010110; // Expected: {'P': 726}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100001; B = 7'b0010110; | Outputs: P=%b | Expected: P=%d",
                 1997,
                 
                 P
                 , 
                 
                 726
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001100; B = 7'b0111010; // Expected: {'P': 696}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001100; B = 7'b0111010; | Outputs: P=%b | Expected: P=%d",
                 1998,
                 
                 P
                 , 
                 
                 696
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101000; B = 7'b1100111; // Expected: {'P': 10712}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101000; B = 7'b1100111; | Outputs: P=%b | Expected: P=%d",
                 1999,
                 
                 P
                 , 
                 
                 10712
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010110; B = 7'b0010000; // Expected: {'P': 1376}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010110; B = 7'b0010000; | Outputs: P=%b | Expected: P=%d",
                 2000,
                 
                 P
                 , 
                 
                 1376
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001011; B = 7'b0001010; // Expected: {'P': 750}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001011; B = 7'b0001010; | Outputs: P=%b | Expected: P=%d",
                 2001,
                 
                 P
                 , 
                 
                 750
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100001; B = 7'b0100111; // Expected: {'P': 3783}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100001; B = 7'b0100111; | Outputs: P=%b | Expected: P=%d",
                 2002,
                 
                 P
                 , 
                 
                 3783
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101010; B = 7'b1011010; // Expected: {'P': 3780}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101010; B = 7'b1011010; | Outputs: P=%b | Expected: P=%d",
                 2003,
                 
                 P
                 , 
                 
                 3780
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011011; B = 7'b1000000; // Expected: {'P': 5824}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011011; B = 7'b1000000; | Outputs: P=%b | Expected: P=%d",
                 2004,
                 
                 P
                 , 
                 
                 5824
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000010; B = 7'b1110110; // Expected: {'P': 236}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000010; B = 7'b1110110; | Outputs: P=%b | Expected: P=%d",
                 2005,
                 
                 P
                 , 
                 
                 236
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111000; B = 7'b1100101; // Expected: {'P': 12120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111000; B = 7'b1100101; | Outputs: P=%b | Expected: P=%d",
                 2006,
                 
                 P
                 , 
                 
                 12120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001110; B = 7'b1100001; // Expected: {'P': 7566}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001110; B = 7'b1100001; | Outputs: P=%b | Expected: P=%d",
                 2007,
                 
                 P
                 , 
                 
                 7566
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100100; B = 7'b0010101; // Expected: {'P': 756}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100100; B = 7'b0010101; | Outputs: P=%b | Expected: P=%d",
                 2008,
                 
                 P
                 , 
                 
                 756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011010; B = 7'b1100110; // Expected: {'P': 2652}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011010; B = 7'b1100110; | Outputs: P=%b | Expected: P=%d",
                 2009,
                 
                 P
                 , 
                 
                 2652
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011010; B = 7'b1100110; // Expected: {'P': 9180}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011010; B = 7'b1100110; | Outputs: P=%b | Expected: P=%d",
                 2010,
                 
                 P
                 , 
                 
                 9180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011000; B = 7'b0000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011000; B = 7'b0000000; | Outputs: P=%b | Expected: P=%d",
                 2011,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110110; B = 7'b0001110; // Expected: {'P': 756}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110110; B = 7'b0001110; | Outputs: P=%b | Expected: P=%d",
                 2012,
                 
                 P
                 , 
                 
                 756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111101; B = 7'b0111110; // Expected: {'P': 7750}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111101; B = 7'b0111110; | Outputs: P=%b | Expected: P=%d",
                 2013,
                 
                 P
                 , 
                 
                 7750
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101010; B = 7'b0001010; // Expected: {'P': 1060}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101010; B = 7'b0001010; | Outputs: P=%b | Expected: P=%d",
                 2014,
                 
                 P
                 , 
                 
                 1060
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110001; B = 7'b1101111; // Expected: {'P': 5439}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110001; B = 7'b1101111; | Outputs: P=%b | Expected: P=%d",
                 2015,
                 
                 P
                 , 
                 
                 5439
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111101; B = 7'b0011011; // Expected: {'P': 1647}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111101; B = 7'b0011011; | Outputs: P=%b | Expected: P=%d",
                 2016,
                 
                 P
                 , 
                 
                 1647
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101111; B = 7'b0101010; // Expected: {'P': 4662}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101111; B = 7'b0101010; | Outputs: P=%b | Expected: P=%d",
                 2017,
                 
                 P
                 , 
                 
                 4662
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001001; B = 7'b1111000; // Expected: {'P': 1080}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001001; B = 7'b1111000; | Outputs: P=%b | Expected: P=%d",
                 2018,
                 
                 P
                 , 
                 
                 1080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101111; B = 7'b0100111; // Expected: {'P': 4329}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101111; B = 7'b0100111; | Outputs: P=%b | Expected: P=%d",
                 2019,
                 
                 P
                 , 
                 
                 4329
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111110; B = 7'b1100101; // Expected: {'P': 12726}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111110; B = 7'b1100101; | Outputs: P=%b | Expected: P=%d",
                 2020,
                 
                 P
                 , 
                 
                 12726
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001001; B = 7'b0110100; // Expected: {'P': 468}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001001; B = 7'b0110100; | Outputs: P=%b | Expected: P=%d",
                 2021,
                 
                 P
                 , 
                 
                 468
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001011; B = 7'b1100111; // Expected: {'P': 7725}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001011; B = 7'b1100111; | Outputs: P=%b | Expected: P=%d",
                 2022,
                 
                 P
                 , 
                 
                 7725
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010001; B = 7'b0010011; // Expected: {'P': 1539}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010001; B = 7'b0010011; | Outputs: P=%b | Expected: P=%d",
                 2023,
                 
                 P
                 , 
                 
                 1539
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100100; B = 7'b0101110; // Expected: {'P': 4600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100100; B = 7'b0101110; | Outputs: P=%b | Expected: P=%d",
                 2024,
                 
                 P
                 , 
                 
                 4600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100100; B = 7'b1111011; // Expected: {'P': 4428}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100100; B = 7'b1111011; | Outputs: P=%b | Expected: P=%d",
                 2025,
                 
                 P
                 , 
                 
                 4428
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011001; B = 7'b1100100; // Expected: {'P': 8900}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011001; B = 7'b1100100; | Outputs: P=%b | Expected: P=%d",
                 2026,
                 
                 P
                 , 
                 
                 8900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010111; B = 7'b0110111; // Expected: {'P': 4785}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010111; B = 7'b0110111; | Outputs: P=%b | Expected: P=%d",
                 2027,
                 
                 P
                 , 
                 
                 4785
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000100; B = 7'b1000011; // Expected: {'P': 4556}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000100; B = 7'b1000011; | Outputs: P=%b | Expected: P=%d",
                 2028,
                 
                 P
                 , 
                 
                 4556
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101101; B = 7'b0001000; // Expected: {'P': 360}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101101; B = 7'b0001000; | Outputs: P=%b | Expected: P=%d",
                 2029,
                 
                 P
                 , 
                 
                 360
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100111; B = 7'b1000100; // Expected: {'P': 7004}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100111; B = 7'b1000100; | Outputs: P=%b | Expected: P=%d",
                 2030,
                 
                 P
                 , 
                 
                 7004
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011010; B = 7'b1001100; // Expected: {'P': 1976}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011010; B = 7'b1001100; | Outputs: P=%b | Expected: P=%d",
                 2031,
                 
                 P
                 , 
                 
                 1976
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101111; B = 7'b0111100; // Expected: {'P': 2820}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101111; B = 7'b0111100; | Outputs: P=%b | Expected: P=%d",
                 2032,
                 
                 P
                 , 
                 
                 2820
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011110; B = 7'b0011110; // Expected: {'P': 2820}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011110; B = 7'b0011110; | Outputs: P=%b | Expected: P=%d",
                 2033,
                 
                 P
                 , 
                 
                 2820
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000011; B = 7'b1010111; // Expected: {'P': 5829}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000011; B = 7'b1010111; | Outputs: P=%b | Expected: P=%d",
                 2034,
                 
                 P
                 , 
                 
                 5829
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000001; B = 7'b0101001; // Expected: {'P': 41}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000001; B = 7'b0101001; | Outputs: P=%b | Expected: P=%d",
                 2035,
                 
                 P
                 , 
                 
                 41
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100101; B = 7'b1111010; // Expected: {'P': 4514}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100101; B = 7'b1111010; | Outputs: P=%b | Expected: P=%d",
                 2036,
                 
                 P
                 , 
                 
                 4514
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011101; B = 7'b1110110; // Expected: {'P': 10974}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011101; B = 7'b1110110; | Outputs: P=%b | Expected: P=%d",
                 2037,
                 
                 P
                 , 
                 
                 10974
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000010; B = 7'b0010111; // Expected: {'P': 1518}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000010; B = 7'b0010111; | Outputs: P=%b | Expected: P=%d",
                 2038,
                 
                 P
                 , 
                 
                 1518
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000110; B = 7'b1101110; // Expected: {'P': 7700}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000110; B = 7'b1101110; | Outputs: P=%b | Expected: P=%d",
                 2039,
                 
                 P
                 , 
                 
                 7700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111111; B = 7'b1111101; // Expected: {'P': 15875}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111111; B = 7'b1111101; | Outputs: P=%b | Expected: P=%d",
                 2040,
                 
                 P
                 , 
                 
                 15875
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001001; B = 7'b1000101; // Expected: {'P': 5037}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001001; B = 7'b1000101; | Outputs: P=%b | Expected: P=%d",
                 2041,
                 
                 P
                 , 
                 
                 5037
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110111; B = 7'b1111001; // Expected: {'P': 14399}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110111; B = 7'b1111001; | Outputs: P=%b | Expected: P=%d",
                 2042,
                 
                 P
                 , 
                 
                 14399
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110010; B = 7'b1101100; // Expected: {'P': 12312}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110010; B = 7'b1101100; | Outputs: P=%b | Expected: P=%d",
                 2043,
                 
                 P
                 , 
                 
                 12312
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110110; B = 7'b0100011; // Expected: {'P': 4130}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110110; B = 7'b0100011; | Outputs: P=%b | Expected: P=%d",
                 2044,
                 
                 P
                 , 
                 
                 4130
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110100; B = 7'b1000001; // Expected: {'P': 3380}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110100; B = 7'b1000001; | Outputs: P=%b | Expected: P=%d",
                 2045,
                 
                 P
                 , 
                 
                 3380
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100110; B = 7'b0000101; // Expected: {'P': 190}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100110; B = 7'b0000101; | Outputs: P=%b | Expected: P=%d",
                 2046,
                 
                 P
                 , 
                 
                 190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100100; B = 7'b0111010; // Expected: {'P': 2088}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100100; B = 7'b0111010; | Outputs: P=%b | Expected: P=%d",
                 2047,
                 
                 P
                 , 
                 
                 2088
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000100; B = 7'b1100000; // Expected: {'P': 384}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000100; B = 7'b1100000; | Outputs: P=%b | Expected: P=%d",
                 2048,
                 
                 P
                 , 
                 
                 384
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111001; B = 7'b0000111; // Expected: {'P': 399}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111001; B = 7'b0000111; | Outputs: P=%b | Expected: P=%d",
                 2049,
                 
                 P
                 , 
                 
                 399
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100100; B = 7'b1010000; // Expected: {'P': 2880}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100100; B = 7'b1010000; | Outputs: P=%b | Expected: P=%d",
                 2050,
                 
                 P
                 , 
                 
                 2880
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000000; B = 7'b1101001; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000000; B = 7'b1101001; | Outputs: P=%b | Expected: P=%d",
                 2051,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010111; B = 7'b0101101; // Expected: {'P': 3915}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010111; B = 7'b0101101; | Outputs: P=%b | Expected: P=%d",
                 2052,
                 
                 P
                 , 
                 
                 3915
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111110; B = 7'b1101001; // Expected: {'P': 13230}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111110; B = 7'b1101001; | Outputs: P=%b | Expected: P=%d",
                 2053,
                 
                 P
                 , 
                 
                 13230
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110110; B = 7'b0010101; // Expected: {'P': 2478}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110110; B = 7'b0010101; | Outputs: P=%b | Expected: P=%d",
                 2054,
                 
                 P
                 , 
                 
                 2478
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110100; B = 7'b1010001; // Expected: {'P': 4212}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110100; B = 7'b1010001; | Outputs: P=%b | Expected: P=%d",
                 2055,
                 
                 P
                 , 
                 
                 4212
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000100; B = 7'b0000001; // Expected: {'P': 68}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000100; B = 7'b0000001; | Outputs: P=%b | Expected: P=%d",
                 2056,
                 
                 P
                 , 
                 
                 68
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101001; B = 7'b0001110; // Expected: {'P': 1470}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101001; B = 7'b0001110; | Outputs: P=%b | Expected: P=%d",
                 2057,
                 
                 P
                 , 
                 
                 1470
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010000; B = 7'b1000000; // Expected: {'P': 5120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010000; B = 7'b1000000; | Outputs: P=%b | Expected: P=%d",
                 2058,
                 
                 P
                 , 
                 
                 5120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011000; B = 7'b0011010; // Expected: {'P': 2288}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011000; B = 7'b0011010; | Outputs: P=%b | Expected: P=%d",
                 2059,
                 
                 P
                 , 
                 
                 2288
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101101; B = 7'b0001011; // Expected: {'P': 1199}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101101; B = 7'b0001011; | Outputs: P=%b | Expected: P=%d",
                 2060,
                 
                 P
                 , 
                 
                 1199
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001100; B = 7'b0011000; // Expected: {'P': 1824}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001100; B = 7'b0011000; | Outputs: P=%b | Expected: P=%d",
                 2061,
                 
                 P
                 , 
                 
                 1824
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001001; B = 7'b0100011; // Expected: {'P': 2555}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001001; B = 7'b0100011; | Outputs: P=%b | Expected: P=%d",
                 2062,
                 
                 P
                 , 
                 
                 2555
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010010; B = 7'b0111111; // Expected: {'P': 5166}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010010; B = 7'b0111111; | Outputs: P=%b | Expected: P=%d",
                 2063,
                 
                 P
                 , 
                 
                 5166
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000111; B = 7'b0000111; // Expected: {'P': 49}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000111; B = 7'b0000111; | Outputs: P=%b | Expected: P=%d",
                 2064,
                 
                 P
                 , 
                 
                 49
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110111; B = 7'b1110101; // Expected: {'P': 6435}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110111; B = 7'b1110101; | Outputs: P=%b | Expected: P=%d",
                 2065,
                 
                 P
                 , 
                 
                 6435
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111001; B = 7'b1000100; // Expected: {'P': 3876}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111001; B = 7'b1000100; | Outputs: P=%b | Expected: P=%d",
                 2066,
                 
                 P
                 , 
                 
                 3876
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010110; B = 7'b0101111; // Expected: {'P': 1034}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010110; B = 7'b0101111; | Outputs: P=%b | Expected: P=%d",
                 2067,
                 
                 P
                 , 
                 
                 1034
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000001; B = 7'b1100001; // Expected: {'P': 97}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000001; B = 7'b1100001; | Outputs: P=%b | Expected: P=%d",
                 2068,
                 
                 P
                 , 
                 
                 97
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110011; B = 7'b0000010; // Expected: {'P': 230}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110011; B = 7'b0000010; | Outputs: P=%b | Expected: P=%d",
                 2069,
                 
                 P
                 , 
                 
                 230
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001000; B = 7'b0011111; // Expected: {'P': 2232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001000; B = 7'b0011111; | Outputs: P=%b | Expected: P=%d",
                 2070,
                 
                 P
                 , 
                 
                 2232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101000; B = 7'b0110110; // Expected: {'P': 5616}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101000; B = 7'b0110110; | Outputs: P=%b | Expected: P=%d",
                 2071,
                 
                 P
                 , 
                 
                 5616
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010110; B = 7'b0010110; // Expected: {'P': 484}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010110; B = 7'b0010110; | Outputs: P=%b | Expected: P=%d",
                 2072,
                 
                 P
                 , 
                 
                 484
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101010; B = 7'b0001110; // Expected: {'P': 1484}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101010; B = 7'b0001110; | Outputs: P=%b | Expected: P=%d",
                 2073,
                 
                 P
                 , 
                 
                 1484
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010000; B = 7'b0000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010000; B = 7'b0000000; | Outputs: P=%b | Expected: P=%d",
                 2074,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100111; B = 7'b1110111; // Expected: {'P': 12257}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100111; B = 7'b1110111; | Outputs: P=%b | Expected: P=%d",
                 2075,
                 
                 P
                 , 
                 
                 12257
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011000; B = 7'b0110101; // Expected: {'P': 4664}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011000; B = 7'b0110101; | Outputs: P=%b | Expected: P=%d",
                 2076,
                 
                 P
                 , 
                 
                 4664
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010001; B = 7'b0100000; // Expected: {'P': 544}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010001; B = 7'b0100000; | Outputs: P=%b | Expected: P=%d",
                 2077,
                 
                 P
                 , 
                 
                 544
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100100; B = 7'b0011100; // Expected: {'P': 1008}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100100; B = 7'b0011100; | Outputs: P=%b | Expected: P=%d",
                 2078,
                 
                 P
                 , 
                 
                 1008
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100001; B = 7'b0111011; // Expected: {'P': 1947}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100001; B = 7'b0111011; | Outputs: P=%b | Expected: P=%d",
                 2079,
                 
                 P
                 , 
                 
                 1947
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110101; B = 7'b0110110; // Expected: {'P': 6318}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110101; B = 7'b0110110; | Outputs: P=%b | Expected: P=%d",
                 2080,
                 
                 P
                 , 
                 
                 6318
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011100; B = 7'b0001001; // Expected: {'P': 828}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011100; B = 7'b0001001; | Outputs: P=%b | Expected: P=%d",
                 2081,
                 
                 P
                 , 
                 
                 828
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000101; B = 7'b1101101; // Expected: {'P': 545}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000101; B = 7'b1101101; | Outputs: P=%b | Expected: P=%d",
                 2082,
                 
                 P
                 , 
                 
                 545
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001100; B = 7'b1010010; // Expected: {'P': 6232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001100; B = 7'b1010010; | Outputs: P=%b | Expected: P=%d",
                 2083,
                 
                 P
                 , 
                 
                 6232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100100; B = 7'b1101111; // Expected: {'P': 3996}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100100; B = 7'b1101111; | Outputs: P=%b | Expected: P=%d",
                 2084,
                 
                 P
                 , 
                 
                 3996
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000110; B = 7'b0101000; // Expected: {'P': 2800}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000110; B = 7'b0101000; | Outputs: P=%b | Expected: P=%d",
                 2085,
                 
                 P
                 , 
                 
                 2800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000100; B = 7'b1011101; // Expected: {'P': 6324}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000100; B = 7'b1011101; | Outputs: P=%b | Expected: P=%d",
                 2086,
                 
                 P
                 , 
                 
                 6324
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000110; B = 7'b0101111; // Expected: {'P': 3290}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000110; B = 7'b0101111; | Outputs: P=%b | Expected: P=%d",
                 2087,
                 
                 P
                 , 
                 
                 3290
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111000; B = 7'b0000100; // Expected: {'P': 480}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111000; B = 7'b0000100; | Outputs: P=%b | Expected: P=%d",
                 2088,
                 
                 P
                 , 
                 
                 480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000101; B = 7'b0011100; // Expected: {'P': 1932}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000101; B = 7'b0011100; | Outputs: P=%b | Expected: P=%d",
                 2089,
                 
                 P
                 , 
                 
                 1932
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110100; B = 7'b0010110; // Expected: {'P': 2552}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110100; B = 7'b0010110; | Outputs: P=%b | Expected: P=%d",
                 2090,
                 
                 P
                 , 
                 
                 2552
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111110; B = 7'b1101000; // Expected: {'P': 6448}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111110; B = 7'b1101000; | Outputs: P=%b | Expected: P=%d",
                 2091,
                 
                 P
                 , 
                 
                 6448
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000110; B = 7'b1111110; // Expected: {'P': 756}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000110; B = 7'b1111110; | Outputs: P=%b | Expected: P=%d",
                 2092,
                 
                 P
                 , 
                 
                 756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000001; B = 7'b1101011; // Expected: {'P': 107}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000001; B = 7'b1101011; | Outputs: P=%b | Expected: P=%d",
                 2093,
                 
                 P
                 , 
                 
                 107
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101001; B = 7'b1101100; // Expected: {'P': 4428}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101001; B = 7'b1101100; | Outputs: P=%b | Expected: P=%d",
                 2094,
                 
                 P
                 , 
                 
                 4428
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001110; B = 7'b0101100; // Expected: {'P': 616}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001110; B = 7'b0101100; | Outputs: P=%b | Expected: P=%d",
                 2095,
                 
                 P
                 , 
                 
                 616
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001011; B = 7'b0110101; // Expected: {'P': 583}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001011; B = 7'b0110101; | Outputs: P=%b | Expected: P=%d",
                 2096,
                 
                 P
                 , 
                 
                 583
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101100; B = 7'b0110101; // Expected: {'P': 2332}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101100; B = 7'b0110101; | Outputs: P=%b | Expected: P=%d",
                 2097,
                 
                 P
                 , 
                 
                 2332
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000101; B = 7'b0000100; // Expected: {'P': 276}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000101; B = 7'b0000100; | Outputs: P=%b | Expected: P=%d",
                 2098,
                 
                 P
                 , 
                 
                 276
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110010; B = 7'b0000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110010; B = 7'b0000000; | Outputs: P=%b | Expected: P=%d",
                 2099,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010011; B = 7'b0101000; // Expected: {'P': 760}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010011; B = 7'b0101000; | Outputs: P=%b | Expected: P=%d",
                 2100,
                 
                 P
                 , 
                 
                 760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101011; B = 7'b1100111; // Expected: {'P': 11021}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101011; B = 7'b1100111; | Outputs: P=%b | Expected: P=%d",
                 2101,
                 
                 P
                 , 
                 
                 11021
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111010; B = 7'b1011110; // Expected: {'P': 5452}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111010; B = 7'b1011110; | Outputs: P=%b | Expected: P=%d",
                 2102,
                 
                 P
                 , 
                 
                 5452
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101111; B = 7'b1000111; // Expected: {'P': 3337}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101111; B = 7'b1000111; | Outputs: P=%b | Expected: P=%d",
                 2103,
                 
                 P
                 , 
                 
                 3337
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001100; B = 7'b0010101; // Expected: {'P': 252}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001100; B = 7'b0010101; | Outputs: P=%b | Expected: P=%d",
                 2104,
                 
                 P
                 , 
                 
                 252
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111111; B = 7'b0111000; // Expected: {'P': 3528}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111111; B = 7'b0111000; | Outputs: P=%b | Expected: P=%d",
                 2105,
                 
                 P
                 , 
                 
                 3528
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100110; B = 7'b0101101; // Expected: {'P': 4590}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100110; B = 7'b0101101; | Outputs: P=%b | Expected: P=%d",
                 2106,
                 
                 P
                 , 
                 
                 4590
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011111; B = 7'b1111111; // Expected: {'P': 12065}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011111; B = 7'b1111111; | Outputs: P=%b | Expected: P=%d",
                 2107,
                 
                 P
                 , 
                 
                 12065
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010000; B = 7'b1010111; // Expected: {'P': 6960}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010000; B = 7'b1010111; | Outputs: P=%b | Expected: P=%d",
                 2108,
                 
                 P
                 , 
                 
                 6960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100110; B = 7'b0011101; // Expected: {'P': 1102}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100110; B = 7'b0011101; | Outputs: P=%b | Expected: P=%d",
                 2109,
                 
                 P
                 , 
                 
                 1102
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110001; B = 7'b0011010; // Expected: {'P': 2938}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110001; B = 7'b0011010; | Outputs: P=%b | Expected: P=%d",
                 2110,
                 
                 P
                 , 
                 
                 2938
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011011; B = 7'b0011010; // Expected: {'P': 2366}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011011; B = 7'b0011010; | Outputs: P=%b | Expected: P=%d",
                 2111,
                 
                 P
                 , 
                 
                 2366
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000110; B = 7'b1011101; // Expected: {'P': 6510}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000110; B = 7'b1011101; | Outputs: P=%b | Expected: P=%d",
                 2112,
                 
                 P
                 , 
                 
                 6510
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011111; B = 7'b0101001; // Expected: {'P': 1271}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011111; B = 7'b0101001; | Outputs: P=%b | Expected: P=%d",
                 2113,
                 
                 P
                 , 
                 
                 1271
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001001; B = 7'b0100100; // Expected: {'P': 2628}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001001; B = 7'b0100100; | Outputs: P=%b | Expected: P=%d",
                 2114,
                 
                 P
                 , 
                 
                 2628
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011110; B = 7'b0101001; // Expected: {'P': 1230}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011110; B = 7'b0101001; | Outputs: P=%b | Expected: P=%d",
                 2115,
                 
                 P
                 , 
                 
                 1230
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100001; B = 7'b0000101; // Expected: {'P': 165}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100001; B = 7'b0000101; | Outputs: P=%b | Expected: P=%d",
                 2116,
                 
                 P
                 , 
                 
                 165
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010011; B = 7'b0110011; // Expected: {'P': 4233}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010011; B = 7'b0110011; | Outputs: P=%b | Expected: P=%d",
                 2117,
                 
                 P
                 , 
                 
                 4233
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111110; B = 7'b1111000; // Expected: {'P': 15120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111110; B = 7'b1111000; | Outputs: P=%b | Expected: P=%d",
                 2118,
                 
                 P
                 , 
                 
                 15120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100100; B = 7'b0001000; // Expected: {'P': 800}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100100; B = 7'b0001000; | Outputs: P=%b | Expected: P=%d",
                 2119,
                 
                 P
                 , 
                 
                 800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001010; B = 7'b1100000; // Expected: {'P': 7104}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001010; B = 7'b1100000; | Outputs: P=%b | Expected: P=%d",
                 2120,
                 
                 P
                 , 
                 
                 7104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110000; B = 7'b0001110; // Expected: {'P': 672}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110000; B = 7'b0001110; | Outputs: P=%b | Expected: P=%d",
                 2121,
                 
                 P
                 , 
                 
                 672
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100000; B = 7'b1001010; // Expected: {'P': 7104}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100000; B = 7'b1001010; | Outputs: P=%b | Expected: P=%d",
                 2122,
                 
                 P
                 , 
                 
                 7104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001000; B = 7'b0111010; // Expected: {'P': 464}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001000; B = 7'b0111010; | Outputs: P=%b | Expected: P=%d",
                 2123,
                 
                 P
                 , 
                 
                 464
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101110; B = 7'b0000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101110; B = 7'b0000000; | Outputs: P=%b | Expected: P=%d",
                 2124,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001011; B = 7'b0011101; // Expected: {'P': 2175}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001011; B = 7'b0011101; | Outputs: P=%b | Expected: P=%d",
                 2125,
                 
                 P
                 , 
                 
                 2175
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001011; B = 7'b1011001; // Expected: {'P': 6675}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001011; B = 7'b1011001; | Outputs: P=%b | Expected: P=%d",
                 2126,
                 
                 P
                 , 
                 
                 6675
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011000; B = 7'b0000110; // Expected: {'P': 144}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011000; B = 7'b0000110; | Outputs: P=%b | Expected: P=%d",
                 2127,
                 
                 P
                 , 
                 
                 144
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111000; B = 7'b1001110; // Expected: {'P': 4368}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111000; B = 7'b1001110; | Outputs: P=%b | Expected: P=%d",
                 2128,
                 
                 P
                 , 
                 
                 4368
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010011; B = 7'b0100010; // Expected: {'P': 2822}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010011; B = 7'b0100010; | Outputs: P=%b | Expected: P=%d",
                 2129,
                 
                 P
                 , 
                 
                 2822
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000000; B = 7'b0011110; // Expected: {'P': 1920}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000000; B = 7'b0011110; | Outputs: P=%b | Expected: P=%d",
                 2130,
                 
                 P
                 , 
                 
                 1920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101000; B = 7'b1111001; // Expected: {'P': 4840}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101000; B = 7'b1111001; | Outputs: P=%b | Expected: P=%d",
                 2131,
                 
                 P
                 , 
                 
                 4840
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100100; B = 7'b0100110; // Expected: {'P': 1368}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100100; B = 7'b0100110; | Outputs: P=%b | Expected: P=%d",
                 2132,
                 
                 P
                 , 
                 
                 1368
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110101; B = 7'b0000011; // Expected: {'P': 351}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110101; B = 7'b0000011; | Outputs: P=%b | Expected: P=%d",
                 2133,
                 
                 P
                 , 
                 
                 351
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010111; B = 7'b0100110; // Expected: {'P': 874}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010111; B = 7'b0100110; | Outputs: P=%b | Expected: P=%d",
                 2134,
                 
                 P
                 , 
                 
                 874
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110010; B = 7'b1001000; // Expected: {'P': 3600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110010; B = 7'b1001000; | Outputs: P=%b | Expected: P=%d",
                 2135,
                 
                 P
                 , 
                 
                 3600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000111; B = 7'b1010101; // Expected: {'P': 595}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000111; B = 7'b1010101; | Outputs: P=%b | Expected: P=%d",
                 2136,
                 
                 P
                 , 
                 
                 595
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001100; B = 7'b1000101; // Expected: {'P': 5244}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001100; B = 7'b1000101; | Outputs: P=%b | Expected: P=%d",
                 2137,
                 
                 P
                 , 
                 
                 5244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110001; B = 7'b0000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110001; B = 7'b0000000; | Outputs: P=%b | Expected: P=%d",
                 2138,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111110; B = 7'b1100010; // Expected: {'P': 12348}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111110; B = 7'b1100010; | Outputs: P=%b | Expected: P=%d",
                 2139,
                 
                 P
                 , 
                 
                 12348
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111110; B = 7'b1010110; // Expected: {'P': 10836}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111110; B = 7'b1010110; | Outputs: P=%b | Expected: P=%d",
                 2140,
                 
                 P
                 , 
                 
                 10836
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111110; B = 7'b1010001; // Expected: {'P': 10206}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111110; B = 7'b1010001; | Outputs: P=%b | Expected: P=%d",
                 2141,
                 
                 P
                 , 
                 
                 10206
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110100; B = 7'b0111100; // Expected: {'P': 3120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110100; B = 7'b0111100; | Outputs: P=%b | Expected: P=%d",
                 2142,
                 
                 P
                 , 
                 
                 3120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111011; B = 7'b1011110; // Expected: {'P': 11562}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111011; B = 7'b1011110; | Outputs: P=%b | Expected: P=%d",
                 2143,
                 
                 P
                 , 
                 
                 11562
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001111; B = 7'b1000011; // Expected: {'P': 1005}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001111; B = 7'b1000011; | Outputs: P=%b | Expected: P=%d",
                 2144,
                 
                 P
                 , 
                 
                 1005
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111010; B = 7'b1101010; // Expected: {'P': 6148}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111010; B = 7'b1101010; | Outputs: P=%b | Expected: P=%d",
                 2145,
                 
                 P
                 , 
                 
                 6148
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011101; B = 7'b0000100; // Expected: {'P': 116}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011101; B = 7'b0000100; | Outputs: P=%b | Expected: P=%d",
                 2146,
                 
                 P
                 , 
                 
                 116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111100; B = 7'b0101101; // Expected: {'P': 5580}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111100; B = 7'b0101101; | Outputs: P=%b | Expected: P=%d",
                 2147,
                 
                 P
                 , 
                 
                 5580
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011111; B = 7'b0111010; // Expected: {'P': 5510}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011111; B = 7'b0111010; | Outputs: P=%b | Expected: P=%d",
                 2148,
                 
                 P
                 , 
                 
                 5510
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011101; B = 7'b0010101; // Expected: {'P': 609}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011101; B = 7'b0010101; | Outputs: P=%b | Expected: P=%d",
                 2149,
                 
                 P
                 , 
                 
                 609
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110010; B = 7'b1101000; // Expected: {'P': 11856}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110010; B = 7'b1101000; | Outputs: P=%b | Expected: P=%d",
                 2150,
                 
                 P
                 , 
                 
                 11856
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111010; B = 7'b0000010; // Expected: {'P': 116}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111010; B = 7'b0000010; | Outputs: P=%b | Expected: P=%d",
                 2151,
                 
                 P
                 , 
                 
                 116
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111011; B = 7'b0101111; // Expected: {'P': 2773}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111011; B = 7'b0101111; | Outputs: P=%b | Expected: P=%d",
                 2152,
                 
                 P
                 , 
                 
                 2773
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111101; B = 7'b1011011; // Expected: {'P': 11375}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111101; B = 7'b1011011; | Outputs: P=%b | Expected: P=%d",
                 2153,
                 
                 P
                 , 
                 
                 11375
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010011; B = 7'b0000101; // Expected: {'P': 95}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010011; B = 7'b0000101; | Outputs: P=%b | Expected: P=%d",
                 2154,
                 
                 P
                 , 
                 
                 95
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101111; B = 7'b0001111; // Expected: {'P': 705}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101111; B = 7'b0001111; | Outputs: P=%b | Expected: P=%d",
                 2155,
                 
                 P
                 , 
                 
                 705
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011111; B = 7'b1001000; // Expected: {'P': 2232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011111; B = 7'b1001000; | Outputs: P=%b | Expected: P=%d",
                 2156,
                 
                 P
                 , 
                 
                 2232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010111; B = 7'b1101110; // Expected: {'P': 2530}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010111; B = 7'b1101110; | Outputs: P=%b | Expected: P=%d",
                 2157,
                 
                 P
                 , 
                 
                 2530
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100011; B = 7'b0111111; // Expected: {'P': 6237}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100011; B = 7'b0111111; | Outputs: P=%b | Expected: P=%d",
                 2158,
                 
                 P
                 , 
                 
                 6237
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010011; B = 7'b1101010; // Expected: {'P': 8798}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010011; B = 7'b1101010; | Outputs: P=%b | Expected: P=%d",
                 2159,
                 
                 P
                 , 
                 
                 8798
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010001; B = 7'b0111110; // Expected: {'P': 1054}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010001; B = 7'b0111110; | Outputs: P=%b | Expected: P=%d",
                 2160,
                 
                 P
                 , 
                 
                 1054
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110001; B = 7'b1000011; // Expected: {'P': 7571}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110001; B = 7'b1000011; | Outputs: P=%b | Expected: P=%d",
                 2161,
                 
                 P
                 , 
                 
                 7571
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101101; B = 7'b0111110; // Expected: {'P': 6758}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101101; B = 7'b0111110; | Outputs: P=%b | Expected: P=%d",
                 2162,
                 
                 P
                 , 
                 
                 6758
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011011; B = 7'b0100100; // Expected: {'P': 972}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011011; B = 7'b0100100; | Outputs: P=%b | Expected: P=%d",
                 2163,
                 
                 P
                 , 
                 
                 972
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011010; B = 7'b0000010; // Expected: {'P': 52}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011010; B = 7'b0000010; | Outputs: P=%b | Expected: P=%d",
                 2164,
                 
                 P
                 , 
                 
                 52
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111101; B = 7'b0110101; // Expected: {'P': 6625}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111101; B = 7'b0110101; | Outputs: P=%b | Expected: P=%d",
                 2165,
                 
                 P
                 , 
                 
                 6625
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001100; B = 7'b1000010; // Expected: {'P': 5016}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001100; B = 7'b1000010; | Outputs: P=%b | Expected: P=%d",
                 2166,
                 
                 P
                 , 
                 
                 5016
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011001; B = 7'b1010000; // Expected: {'P': 2000}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011001; B = 7'b1010000; | Outputs: P=%b | Expected: P=%d",
                 2167,
                 
                 P
                 , 
                 
                 2000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001000; B = 7'b0111100; // Expected: {'P': 4320}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001000; B = 7'b0111100; | Outputs: P=%b | Expected: P=%d",
                 2168,
                 
                 P
                 , 
                 
                 4320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100011; B = 7'b0111000; // Expected: {'P': 1960}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100011; B = 7'b0111000; | Outputs: P=%b | Expected: P=%d",
                 2169,
                 
                 P
                 , 
                 
                 1960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000000; B = 7'b0001100; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000000; B = 7'b0001100; | Outputs: P=%b | Expected: P=%d",
                 2170,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010010; B = 7'b0100100; // Expected: {'P': 2952}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010010; B = 7'b0100100; | Outputs: P=%b | Expected: P=%d",
                 2171,
                 
                 P
                 , 
                 
                 2952
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110011; B = 7'b1001110; // Expected: {'P': 8970}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110011; B = 7'b1001110; | Outputs: P=%b | Expected: P=%d",
                 2172,
                 
                 P
                 , 
                 
                 8970
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100000; B = 7'b1010101; // Expected: {'P': 2720}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100000; B = 7'b1010101; | Outputs: P=%b | Expected: P=%d",
                 2173,
                 
                 P
                 , 
                 
                 2720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001011; B = 7'b1110110; // Expected: {'P': 8850}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001011; B = 7'b1110110; | Outputs: P=%b | Expected: P=%d",
                 2174,
                 
                 P
                 , 
                 
                 8850
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010101; B = 7'b0000010; // Expected: {'P': 170}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010101; B = 7'b0000010; | Outputs: P=%b | Expected: P=%d",
                 2175,
                 
                 P
                 , 
                 
                 170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110010; B = 7'b1100110; // Expected: {'P': 5100}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110010; B = 7'b1100110; | Outputs: P=%b | Expected: P=%d",
                 2176,
                 
                 P
                 , 
                 
                 5100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110100; B = 7'b1011010; // Expected: {'P': 10440}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110100; B = 7'b1011010; | Outputs: P=%b | Expected: P=%d",
                 2177,
                 
                 P
                 , 
                 
                 10440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000101; B = 7'b0101100; // Expected: {'P': 3036}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000101; B = 7'b0101100; | Outputs: P=%b | Expected: P=%d",
                 2178,
                 
                 P
                 , 
                 
                 3036
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111100; B = 7'b0000001; // Expected: {'P': 124}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111100; B = 7'b0000001; | Outputs: P=%b | Expected: P=%d",
                 2179,
                 
                 P
                 , 
                 
                 124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010000; B = 7'b0110100; // Expected: {'P': 4160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010000; B = 7'b0110100; | Outputs: P=%b | Expected: P=%d",
                 2180,
                 
                 P
                 , 
                 
                 4160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010101; B = 7'b1010001; // Expected: {'P': 6885}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010101; B = 7'b1010001; | Outputs: P=%b | Expected: P=%d",
                 2181,
                 
                 P
                 , 
                 
                 6885
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101101; B = 7'b0100100; // Expected: {'P': 1620}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101101; B = 7'b0100100; | Outputs: P=%b | Expected: P=%d",
                 2182,
                 
                 P
                 , 
                 
                 1620
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110101; B = 7'b1101101; // Expected: {'P': 5777}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110101; B = 7'b1101101; | Outputs: P=%b | Expected: P=%d",
                 2183,
                 
                 P
                 , 
                 
                 5777
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110010; B = 7'b1100010; // Expected: {'P': 4900}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110010; B = 7'b1100010; | Outputs: P=%b | Expected: P=%d",
                 2184,
                 
                 P
                 , 
                 
                 4900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000100; B = 7'b1010000; // Expected: {'P': 5440}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000100; B = 7'b1010000; | Outputs: P=%b | Expected: P=%d",
                 2185,
                 
                 P
                 , 
                 
                 5440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111101; B = 7'b0101111; // Expected: {'P': 2867}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111101; B = 7'b0101111; | Outputs: P=%b | Expected: P=%d",
                 2186,
                 
                 P
                 , 
                 
                 2867
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001111; B = 7'b0100111; // Expected: {'P': 3081}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001111; B = 7'b0100111; | Outputs: P=%b | Expected: P=%d",
                 2187,
                 
                 P
                 , 
                 
                 3081
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011111; B = 7'b1010110; // Expected: {'P': 8170}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011111; B = 7'b1010110; | Outputs: P=%b | Expected: P=%d",
                 2188,
                 
                 P
                 , 
                 
                 8170
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110011; B = 7'b1001010; // Expected: {'P': 8510}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110011; B = 7'b1001010; | Outputs: P=%b | Expected: P=%d",
                 2189,
                 
                 P
                 , 
                 
                 8510
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110110; B = 7'b0011000; // Expected: {'P': 1296}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110110; B = 7'b0011000; | Outputs: P=%b | Expected: P=%d",
                 2190,
                 
                 P
                 , 
                 
                 1296
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111011; B = 7'b0011111; // Expected: {'P': 3813}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111011; B = 7'b0011111; | Outputs: P=%b | Expected: P=%d",
                 2191,
                 
                 P
                 , 
                 
                 3813
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011100; B = 7'b0101000; // Expected: {'P': 1120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011100; B = 7'b0101000; | Outputs: P=%b | Expected: P=%d",
                 2192,
                 
                 P
                 , 
                 
                 1120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001101; B = 7'b0100010; // Expected: {'P': 2618}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001101; B = 7'b0100010; | Outputs: P=%b | Expected: P=%d",
                 2193,
                 
                 P
                 , 
                 
                 2618
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000000; B = 7'b1110001; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000000; B = 7'b1110001; | Outputs: P=%b | Expected: P=%d",
                 2194,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000000; B = 7'b1011001; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000000; B = 7'b1011001; | Outputs: P=%b | Expected: P=%d",
                 2195,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100101; B = 7'b0011000; // Expected: {'P': 888}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100101; B = 7'b0011000; | Outputs: P=%b | Expected: P=%d",
                 2196,
                 
                 P
                 , 
                 
                 888
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000101; B = 7'b0100110; // Expected: {'P': 2622}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000101; B = 7'b0100110; | Outputs: P=%b | Expected: P=%d",
                 2197,
                 
                 P
                 , 
                 
                 2622
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000001; B = 7'b1000101; // Expected: {'P': 69}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000001; B = 7'b1000101; | Outputs: P=%b | Expected: P=%d",
                 2198,
                 
                 P
                 , 
                 
                 69
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011011; B = 7'b1110110; // Expected: {'P': 10738}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011011; B = 7'b1110110; | Outputs: P=%b | Expected: P=%d",
                 2199,
                 
                 P
                 , 
                 
                 10738
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011000; B = 7'b0110111; // Expected: {'P': 1320}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011000; B = 7'b0110111; | Outputs: P=%b | Expected: P=%d",
                 2200,
                 
                 P
                 , 
                 
                 1320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111000; B = 7'b1101101; // Expected: {'P': 6104}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111000; B = 7'b1101101; | Outputs: P=%b | Expected: P=%d",
                 2201,
                 
                 P
                 , 
                 
                 6104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011100; B = 7'b1111111; // Expected: {'P': 3556}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011100; B = 7'b1111111; | Outputs: P=%b | Expected: P=%d",
                 2202,
                 
                 P
                 , 
                 
                 3556
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111110; B = 7'b0000101; // Expected: {'P': 310}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111110; B = 7'b0000101; | Outputs: P=%b | Expected: P=%d",
                 2203,
                 
                 P
                 , 
                 
                 310
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100001; B = 7'b1111001; // Expected: {'P': 11737}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100001; B = 7'b1111001; | Outputs: P=%b | Expected: P=%d",
                 2204,
                 
                 P
                 , 
                 
                 11737
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000110; B = 7'b0110011; // Expected: {'P': 306}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000110; B = 7'b0110011; | Outputs: P=%b | Expected: P=%d",
                 2205,
                 
                 P
                 , 
                 
                 306
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000111; B = 7'b1001100; // Expected: {'P': 532}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000111; B = 7'b1001100; | Outputs: P=%b | Expected: P=%d",
                 2206,
                 
                 P
                 , 
                 
                 532
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010000; B = 7'b1101011; // Expected: {'P': 1712}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010000; B = 7'b1101011; | Outputs: P=%b | Expected: P=%d",
                 2207,
                 
                 P
                 , 
                 
                 1712
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010101; B = 7'b1011111; // Expected: {'P': 1995}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010101; B = 7'b1011111; | Outputs: P=%b | Expected: P=%d",
                 2208,
                 
                 P
                 , 
                 
                 1995
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110101; B = 7'b1110101; // Expected: {'P': 13689}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110101; B = 7'b1110101; | Outputs: P=%b | Expected: P=%d",
                 2209,
                 
                 P
                 , 
                 
                 13689
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001011; B = 7'b0000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001011; B = 7'b0000000; | Outputs: P=%b | Expected: P=%d",
                 2210,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110010; B = 7'b1010100; // Expected: {'P': 9576}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110010; B = 7'b1010100; | Outputs: P=%b | Expected: P=%d",
                 2211,
                 
                 P
                 , 
                 
                 9576
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011010; B = 7'b1011000; // Expected: {'P': 7920}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011010; B = 7'b1011000; | Outputs: P=%b | Expected: P=%d",
                 2212,
                 
                 P
                 , 
                 
                 7920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011010; B = 7'b1010111; // Expected: {'P': 2262}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011010; B = 7'b1010111; | Outputs: P=%b | Expected: P=%d",
                 2213,
                 
                 P
                 , 
                 
                 2262
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010100; B = 7'b0101101; // Expected: {'P': 900}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010100; B = 7'b0101101; | Outputs: P=%b | Expected: P=%d",
                 2214,
                 
                 P
                 , 
                 
                 900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011100; B = 7'b0011000; // Expected: {'P': 672}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011100; B = 7'b0011000; | Outputs: P=%b | Expected: P=%d",
                 2215,
                 
                 P
                 , 
                 
                 672
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110000; B = 7'b1000100; // Expected: {'P': 3264}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110000; B = 7'b1000100; | Outputs: P=%b | Expected: P=%d",
                 2216,
                 
                 P
                 , 
                 
                 3264
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101001; B = 7'b1100111; // Expected: {'P': 10815}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101001; B = 7'b1100111; | Outputs: P=%b | Expected: P=%d",
                 2217,
                 
                 P
                 , 
                 
                 10815
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111101; B = 7'b0100000; // Expected: {'P': 4000}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111101; B = 7'b0100000; | Outputs: P=%b | Expected: P=%d",
                 2218,
                 
                 P
                 , 
                 
                 4000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101010; B = 7'b1010100; // Expected: {'P': 3528}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101010; B = 7'b1010100; | Outputs: P=%b | Expected: P=%d",
                 2219,
                 
                 P
                 , 
                 
                 3528
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010000; B = 7'b1010100; // Expected: {'P': 1344}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010000; B = 7'b1010100; | Outputs: P=%b | Expected: P=%d",
                 2220,
                 
                 P
                 , 
                 
                 1344
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010110; B = 7'b0100101; // Expected: {'P': 3182}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010110; B = 7'b0100101; | Outputs: P=%b | Expected: P=%d",
                 2221,
                 
                 P
                 , 
                 
                 3182
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101100; B = 7'b0011110; // Expected: {'P': 1320}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101100; B = 7'b0011110; | Outputs: P=%b | Expected: P=%d",
                 2222,
                 
                 P
                 , 
                 
                 1320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000001; B = 7'b0101110; // Expected: {'P': 46}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000001; B = 7'b0101110; | Outputs: P=%b | Expected: P=%d",
                 2223,
                 
                 P
                 , 
                 
                 46
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001101; B = 7'b1111011; // Expected: {'P': 1599}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001101; B = 7'b1111011; | Outputs: P=%b | Expected: P=%d",
                 2224,
                 
                 P
                 , 
                 
                 1599
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110101; B = 7'b0100010; // Expected: {'P': 3978}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110101; B = 7'b0100010; | Outputs: P=%b | Expected: P=%d",
                 2225,
                 
                 P
                 , 
                 
                 3978
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101011; B = 7'b0001000; // Expected: {'P': 344}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101011; B = 7'b0001000; | Outputs: P=%b | Expected: P=%d",
                 2226,
                 
                 P
                 , 
                 
                 344
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011110; B = 7'b0011011; // Expected: {'P': 2538}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011110; B = 7'b0011011; | Outputs: P=%b | Expected: P=%d",
                 2227,
                 
                 P
                 , 
                 
                 2538
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001111; B = 7'b0000011; // Expected: {'P': 45}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001111; B = 7'b0000011; | Outputs: P=%b | Expected: P=%d",
                 2228,
                 
                 P
                 , 
                 
                 45
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111010; B = 7'b0000011; // Expected: {'P': 174}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111010; B = 7'b0000011; | Outputs: P=%b | Expected: P=%d",
                 2229,
                 
                 P
                 , 
                 
                 174
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110011; B = 7'b1010011; // Expected: {'P': 4233}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110011; B = 7'b1010011; | Outputs: P=%b | Expected: P=%d",
                 2230,
                 
                 P
                 , 
                 
                 4233
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100111; B = 7'b1111101; // Expected: {'P': 4875}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100111; B = 7'b1111101; | Outputs: P=%b | Expected: P=%d",
                 2231,
                 
                 P
                 , 
                 
                 4875
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100000; B = 7'b1011100; // Expected: {'P': 2944}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100000; B = 7'b1011100; | Outputs: P=%b | Expected: P=%d",
                 2232,
                 
                 P
                 , 
                 
                 2944
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101100; B = 7'b0000001; // Expected: {'P': 44}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101100; B = 7'b0000001; | Outputs: P=%b | Expected: P=%d",
                 2233,
                 
                 P
                 , 
                 
                 44
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101000; B = 7'b1100111; // Expected: {'P': 4120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101000; B = 7'b1100111; | Outputs: P=%b | Expected: P=%d",
                 2234,
                 
                 P
                 , 
                 
                 4120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010101; B = 7'b0101101; // Expected: {'P': 3825}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010101; B = 7'b0101101; | Outputs: P=%b | Expected: P=%d",
                 2235,
                 
                 P
                 , 
                 
                 3825
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011000; B = 7'b0001001; // Expected: {'P': 792}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011000; B = 7'b0001001; | Outputs: P=%b | Expected: P=%d",
                 2236,
                 
                 P
                 , 
                 
                 792
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011111; B = 7'b1100100; // Expected: {'P': 9500}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011111; B = 7'b1100100; | Outputs: P=%b | Expected: P=%d",
                 2237,
                 
                 P
                 , 
                 
                 9500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010010; B = 7'b0010011; // Expected: {'P': 342}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010010; B = 7'b0010011; | Outputs: P=%b | Expected: P=%d",
                 2238,
                 
                 P
                 , 
                 
                 342
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101111; B = 7'b1111100; // Expected: {'P': 5828}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101111; B = 7'b1111100; | Outputs: P=%b | Expected: P=%d",
                 2239,
                 
                 P
                 , 
                 
                 5828
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010111; B = 7'b0011111; // Expected: {'P': 713}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010111; B = 7'b0011111; | Outputs: P=%b | Expected: P=%d",
                 2240,
                 
                 P
                 , 
                 
                 713
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111001; B = 7'b1110100; // Expected: {'P': 14036}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111001; B = 7'b1110100; | Outputs: P=%b | Expected: P=%d",
                 2241,
                 
                 P
                 , 
                 
                 14036
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100111; B = 7'b0001010; // Expected: {'P': 1030}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100111; B = 7'b0001010; | Outputs: P=%b | Expected: P=%d",
                 2242,
                 
                 P
                 , 
                 
                 1030
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101111; B = 7'b0100000; // Expected: {'P': 1504}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101111; B = 7'b0100000; | Outputs: P=%b | Expected: P=%d",
                 2243,
                 
                 P
                 , 
                 
                 1504
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010000; B = 7'b1000011; // Expected: {'P': 1072}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010000; B = 7'b1000011; | Outputs: P=%b | Expected: P=%d",
                 2244,
                 
                 P
                 , 
                 
                 1072
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010100; B = 7'b0011001; // Expected: {'P': 2100}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010100; B = 7'b0011001; | Outputs: P=%b | Expected: P=%d",
                 2245,
                 
                 P
                 , 
                 
                 2100
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011010; B = 7'b0010110; // Expected: {'P': 1980}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011010; B = 7'b0010110; | Outputs: P=%b | Expected: P=%d",
                 2246,
                 
                 P
                 , 
                 
                 1980
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111001; B = 7'b1111011; // Expected: {'P': 14883}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111001; B = 7'b1111011; | Outputs: P=%b | Expected: P=%d",
                 2247,
                 
                 P
                 , 
                 
                 14883
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101110; B = 7'b1001111; // Expected: {'P': 8690}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101110; B = 7'b1001111; | Outputs: P=%b | Expected: P=%d",
                 2248,
                 
                 P
                 , 
                 
                 8690
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011001; B = 7'b1011111; // Expected: {'P': 2375}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011001; B = 7'b1011111; | Outputs: P=%b | Expected: P=%d",
                 2249,
                 
                 P
                 , 
                 
                 2375
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100011; B = 7'b0000110; // Expected: {'P': 210}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100011; B = 7'b0000110; | Outputs: P=%b | Expected: P=%d",
                 2250,
                 
                 P
                 , 
                 
                 210
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110111; B = 7'b0000110; // Expected: {'P': 714}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110111; B = 7'b0000110; | Outputs: P=%b | Expected: P=%d",
                 2251,
                 
                 P
                 , 
                 
                 714
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111111; B = 7'b0001100; // Expected: {'P': 756}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111111; B = 7'b0001100; | Outputs: P=%b | Expected: P=%d",
                 2252,
                 
                 P
                 , 
                 
                 756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000101; B = 7'b0000101; // Expected: {'P': 345}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000101; B = 7'b0000101; | Outputs: P=%b | Expected: P=%d",
                 2253,
                 
                 P
                 , 
                 
                 345
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000111; B = 7'b1011010; // Expected: {'P': 6390}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000111; B = 7'b1011010; | Outputs: P=%b | Expected: P=%d",
                 2254,
                 
                 P
                 , 
                 
                 6390
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001010; B = 7'b1001111; // Expected: {'P': 5846}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001010; B = 7'b1001111; | Outputs: P=%b | Expected: P=%d",
                 2255,
                 
                 P
                 , 
                 
                 5846
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011110; B = 7'b1001000; // Expected: {'P': 2160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011110; B = 7'b1001000; | Outputs: P=%b | Expected: P=%d",
                 2256,
                 
                 P
                 , 
                 
                 2160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000110; B = 7'b1011111; // Expected: {'P': 6650}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000110; B = 7'b1011111; | Outputs: P=%b | Expected: P=%d",
                 2257,
                 
                 P
                 , 
                 
                 6650
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101011; B = 7'b0000001; // Expected: {'P': 43}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101011; B = 7'b0000001; | Outputs: P=%b | Expected: P=%d",
                 2258,
                 
                 P
                 , 
                 
                 43
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100000; B = 7'b1110110; // Expected: {'P': 3776}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100000; B = 7'b1110110; | Outputs: P=%b | Expected: P=%d",
                 2259,
                 
                 P
                 , 
                 
                 3776
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000101; B = 7'b0010010; // Expected: {'P': 90}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000101; B = 7'b0010010; | Outputs: P=%b | Expected: P=%d",
                 2260,
                 
                 P
                 , 
                 
                 90
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011000; B = 7'b0101111; // Expected: {'P': 1128}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011000; B = 7'b0101111; | Outputs: P=%b | Expected: P=%d",
                 2261,
                 
                 P
                 , 
                 
                 1128
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011101; B = 7'b0110010; // Expected: {'P': 4650}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011101; B = 7'b0110010; | Outputs: P=%b | Expected: P=%d",
                 2262,
                 
                 P
                 , 
                 
                 4650
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000010; B = 7'b1001101; // Expected: {'P': 5082}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000010; B = 7'b1001101; | Outputs: P=%b | Expected: P=%d",
                 2263,
                 
                 P
                 , 
                 
                 5082
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111001; B = 7'b0000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111001; B = 7'b0000000; | Outputs: P=%b | Expected: P=%d",
                 2264,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000110; B = 7'b1111111; // Expected: {'P': 762}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000110; B = 7'b1111111; | Outputs: P=%b | Expected: P=%d",
                 2265,
                 
                 P
                 , 
                 
                 762
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110000; B = 7'b0101111; // Expected: {'P': 2256}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110000; B = 7'b0101111; | Outputs: P=%b | Expected: P=%d",
                 2266,
                 
                 P
                 , 
                 
                 2256
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001100; B = 7'b1111111; // Expected: {'P': 1524}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001100; B = 7'b1111111; | Outputs: P=%b | Expected: P=%d",
                 2267,
                 
                 P
                 , 
                 
                 1524
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101111; B = 7'b0110100; // Expected: {'P': 5772}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101111; B = 7'b0110100; | Outputs: P=%b | Expected: P=%d",
                 2268,
                 
                 P
                 , 
                 
                 5772
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100011; B = 7'b1111001; // Expected: {'P': 11979}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100011; B = 7'b1111001; | Outputs: P=%b | Expected: P=%d",
                 2269,
                 
                 P
                 , 
                 
                 11979
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111001; B = 7'b0011111; // Expected: {'P': 3751}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111001; B = 7'b0011111; | Outputs: P=%b | Expected: P=%d",
                 2270,
                 
                 P
                 , 
                 
                 3751
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001001; B = 7'b1011101; // Expected: {'P': 6789}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001001; B = 7'b1011101; | Outputs: P=%b | Expected: P=%d",
                 2271,
                 
                 P
                 , 
                 
                 6789
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100000; B = 7'b0001100; // Expected: {'P': 1152}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100000; B = 7'b0001100; | Outputs: P=%b | Expected: P=%d",
                 2272,
                 
                 P
                 , 
                 
                 1152
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111010; B = 7'b0101011; // Expected: {'P': 5246}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111010; B = 7'b0101011; | Outputs: P=%b | Expected: P=%d",
                 2273,
                 
                 P
                 , 
                 
                 5246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000011; B = 7'b1001111; // Expected: {'P': 237}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000011; B = 7'b1001111; | Outputs: P=%b | Expected: P=%d",
                 2274,
                 
                 P
                 , 
                 
                 237
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001101; B = 7'b0111001; // Expected: {'P': 4389}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001101; B = 7'b0111001; | Outputs: P=%b | Expected: P=%d",
                 2275,
                 
                 P
                 , 
                 
                 4389
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010110; B = 7'b1101001; // Expected: {'P': 9030}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010110; B = 7'b1101001; | Outputs: P=%b | Expected: P=%d",
                 2276,
                 
                 P
                 , 
                 
                 9030
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110010; B = 7'b1010111; // Expected: {'P': 9918}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110010; B = 7'b1010111; | Outputs: P=%b | Expected: P=%d",
                 2277,
                 
                 P
                 , 
                 
                 9918
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111011; B = 7'b0111101; // Expected: {'P': 7503}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111011; B = 7'b0111101; | Outputs: P=%b | Expected: P=%d",
                 2278,
                 
                 P
                 , 
                 
                 7503
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010010; B = 7'b0111011; // Expected: {'P': 4838}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010010; B = 7'b0111011; | Outputs: P=%b | Expected: P=%d",
                 2279,
                 
                 P
                 , 
                 
                 4838
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111011; B = 7'b0011011; // Expected: {'P': 1593}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111011; B = 7'b0011011; | Outputs: P=%b | Expected: P=%d",
                 2280,
                 
                 P
                 , 
                 
                 1593
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111111; B = 7'b0001110; // Expected: {'P': 882}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111111; B = 7'b0001110; | Outputs: P=%b | Expected: P=%d",
                 2281,
                 
                 P
                 , 
                 
                 882
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110110; B = 7'b1100001; // Expected: {'P': 5238}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110110; B = 7'b1100001; | Outputs: P=%b | Expected: P=%d",
                 2282,
                 
                 P
                 , 
                 
                 5238
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100110; B = 7'b0100101; // Expected: {'P': 3774}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100110; B = 7'b0100101; | Outputs: P=%b | Expected: P=%d",
                 2283,
                 
                 P
                 , 
                 
                 3774
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000011; B = 7'b1110011; // Expected: {'P': 345}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000011; B = 7'b1110011; | Outputs: P=%b | Expected: P=%d",
                 2284,
                 
                 P
                 , 
                 
                 345
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101100; B = 7'b1111111; // Expected: {'P': 13716}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101100; B = 7'b1111111; | Outputs: P=%b | Expected: P=%d",
                 2285,
                 
                 P
                 , 
                 
                 13716
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000010; B = 7'b0000001; // Expected: {'P': 66}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000010; B = 7'b0000001; | Outputs: P=%b | Expected: P=%d",
                 2286,
                 
                 P
                 , 
                 
                 66
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111010; B = 7'b0101010; // Expected: {'P': 5124}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111010; B = 7'b0101010; | Outputs: P=%b | Expected: P=%d",
                 2287,
                 
                 P
                 , 
                 
                 5124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010010; B = 7'b0001000; // Expected: {'P': 656}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010010; B = 7'b0001000; | Outputs: P=%b | Expected: P=%d",
                 2288,
                 
                 P
                 , 
                 
                 656
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111000; B = 7'b0101100; // Expected: {'P': 5280}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111000; B = 7'b0101100; | Outputs: P=%b | Expected: P=%d",
                 2289,
                 
                 P
                 , 
                 
                 5280
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000000; B = 7'b0111001; // Expected: {'P': 3648}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000000; B = 7'b0111001; | Outputs: P=%b | Expected: P=%d",
                 2290,
                 
                 P
                 , 
                 
                 3648
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011011; B = 7'b1101001; // Expected: {'P': 9555}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011011; B = 7'b1101001; | Outputs: P=%b | Expected: P=%d",
                 2291,
                 
                 P
                 , 
                 
                 9555
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111010; B = 7'b1101000; // Expected: {'P': 6032}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111010; B = 7'b1101000; | Outputs: P=%b | Expected: P=%d",
                 2292,
                 
                 P
                 , 
                 
                 6032
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111110; B = 7'b0101010; // Expected: {'P': 2604}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111110; B = 7'b0101010; | Outputs: P=%b | Expected: P=%d",
                 2293,
                 
                 P
                 , 
                 
                 2604
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111001; B = 7'b1011101; // Expected: {'P': 11253}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111001; B = 7'b1011101; | Outputs: P=%b | Expected: P=%d",
                 2294,
                 
                 P
                 , 
                 
                 11253
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101001; B = 7'b1000100; // Expected: {'P': 7140}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101001; B = 7'b1000100; | Outputs: P=%b | Expected: P=%d",
                 2295,
                 
                 P
                 , 
                 
                 7140
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011110; B = 7'b1110000; // Expected: {'P': 10528}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011110; B = 7'b1110000; | Outputs: P=%b | Expected: P=%d",
                 2296,
                 
                 P
                 , 
                 
                 10528
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001101; B = 7'b0000001; // Expected: {'P': 77}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001101; B = 7'b0000001; | Outputs: P=%b | Expected: P=%d",
                 2297,
                 
                 P
                 , 
                 
                 77
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010111; B = 7'b1111001; // Expected: {'P': 10527}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010111; B = 7'b1111001; | Outputs: P=%b | Expected: P=%d",
                 2298,
                 
                 P
                 , 
                 
                 10527
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011111; B = 7'b1001111; // Expected: {'P': 7505}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011111; B = 7'b1001111; | Outputs: P=%b | Expected: P=%d",
                 2299,
                 
                 P
                 , 
                 
                 7505
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100001; B = 7'b0000001; // Expected: {'P': 33}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100001; B = 7'b0000001; | Outputs: P=%b | Expected: P=%d",
                 2300,
                 
                 P
                 , 
                 
                 33
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101000; B = 7'b0101100; // Expected: {'P': 4576}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101000; B = 7'b0101100; | Outputs: P=%b | Expected: P=%d",
                 2301,
                 
                 P
                 , 
                 
                 4576
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001000; B = 7'b0100110; // Expected: {'P': 304}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001000; B = 7'b0100110; | Outputs: P=%b | Expected: P=%d",
                 2302,
                 
                 P
                 , 
                 
                 304
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001000; B = 7'b1000110; // Expected: {'P': 560}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001000; B = 7'b1000110; | Outputs: P=%b | Expected: P=%d",
                 2303,
                 
                 P
                 , 
                 
                 560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001001; B = 7'b1111101; // Expected: {'P': 1125}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001001; B = 7'b1111101; | Outputs: P=%b | Expected: P=%d",
                 2304,
                 
                 P
                 , 
                 
                 1125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010110; B = 7'b1010000; // Expected: {'P': 1760}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010110; B = 7'b1010000; | Outputs: P=%b | Expected: P=%d",
                 2305,
                 
                 P
                 , 
                 
                 1760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101100; B = 7'b0101010; // Expected: {'P': 4536}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101100; B = 7'b0101010; | Outputs: P=%b | Expected: P=%d",
                 2306,
                 
                 P
                 , 
                 
                 4536
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011010; B = 7'b1011010; // Expected: {'P': 2340}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011010; B = 7'b1011010; | Outputs: P=%b | Expected: P=%d",
                 2307,
                 
                 P
                 , 
                 
                 2340
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100000; B = 7'b0100100; // Expected: {'P': 3456}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100000; B = 7'b0100100; | Outputs: P=%b | Expected: P=%d",
                 2308,
                 
                 P
                 , 
                 
                 3456
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011110; B = 7'b0110000; // Expected: {'P': 1440}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011110; B = 7'b0110000; | Outputs: P=%b | Expected: P=%d",
                 2309,
                 
                 P
                 , 
                 
                 1440
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111000; B = 7'b0101101; // Expected: {'P': 5400}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111000; B = 7'b0101101; | Outputs: P=%b | Expected: P=%d",
                 2310,
                 
                 P
                 , 
                 
                 5400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000011; B = 7'b1001101; // Expected: {'P': 231}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000011; B = 7'b1001101; | Outputs: P=%b | Expected: P=%d",
                 2311,
                 
                 P
                 , 
                 
                 231
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100101; B = 7'b0000110; // Expected: {'P': 222}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100101; B = 7'b0000110; | Outputs: P=%b | Expected: P=%d",
                 2312,
                 
                 P
                 , 
                 
                 222
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010011; B = 7'b0100110; // Expected: {'P': 3154}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010011; B = 7'b0100110; | Outputs: P=%b | Expected: P=%d",
                 2313,
                 
                 P
                 , 
                 
                 3154
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110001; B = 7'b0010111; // Expected: {'P': 1127}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110001; B = 7'b0010111; | Outputs: P=%b | Expected: P=%d",
                 2314,
                 
                 P
                 , 
                 
                 1127
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111001; B = 7'b0001110; // Expected: {'P': 1694}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111001; B = 7'b0001110; | Outputs: P=%b | Expected: P=%d",
                 2315,
                 
                 P
                 , 
                 
                 1694
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010100; B = 7'b1010111; // Expected: {'P': 7308}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010100; B = 7'b1010111; | Outputs: P=%b | Expected: P=%d",
                 2316,
                 
                 P
                 , 
                 
                 7308
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011000; B = 7'b1100000; // Expected: {'P': 2304}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011000; B = 7'b1100000; | Outputs: P=%b | Expected: P=%d",
                 2317,
                 
                 P
                 , 
                 
                 2304
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110101; B = 7'b0000110; // Expected: {'P': 702}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110101; B = 7'b0000110; | Outputs: P=%b | Expected: P=%d",
                 2318,
                 
                 P
                 , 
                 
                 702
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100111; B = 7'b0000101; // Expected: {'P': 515}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100111; B = 7'b0000101; | Outputs: P=%b | Expected: P=%d",
                 2319,
                 
                 P
                 , 
                 
                 515
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001001; B = 7'b1011010; // Expected: {'P': 6570}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001001; B = 7'b1011010; | Outputs: P=%b | Expected: P=%d",
                 2320,
                 
                 P
                 , 
                 
                 6570
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111111; B = 7'b0111101; // Expected: {'P': 3843}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111111; B = 7'b0111101; | Outputs: P=%b | Expected: P=%d",
                 2321,
                 
                 P
                 , 
                 
                 3843
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000010; B = 7'b1011010; // Expected: {'P': 180}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000010; B = 7'b1011010; | Outputs: P=%b | Expected: P=%d",
                 2322,
                 
                 P
                 , 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000110; B = 7'b1110001; // Expected: {'P': 7910}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000110; B = 7'b1110001; | Outputs: P=%b | Expected: P=%d",
                 2323,
                 
                 P
                 , 
                 
                 7910
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001011; B = 7'b1001011; // Expected: {'P': 5625}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001011; B = 7'b1001011; | Outputs: P=%b | Expected: P=%d",
                 2324,
                 
                 P
                 , 
                 
                 5625
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110100; B = 7'b1011100; // Expected: {'P': 10672}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110100; B = 7'b1011100; | Outputs: P=%b | Expected: P=%d",
                 2325,
                 
                 P
                 , 
                 
                 10672
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101101; B = 7'b1111100; // Expected: {'P': 13516}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101101; B = 7'b1111100; | Outputs: P=%b | Expected: P=%d",
                 2326,
                 
                 P
                 , 
                 
                 13516
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000001; B = 7'b1000111; // Expected: {'P': 4615}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000001; B = 7'b1000111; | Outputs: P=%b | Expected: P=%d",
                 2327,
                 
                 P
                 , 
                 
                 4615
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000111; B = 7'b1100110; // Expected: {'P': 714}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000111; B = 7'b1100110; | Outputs: P=%b | Expected: P=%d",
                 2328,
                 
                 P
                 , 
                 
                 714
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000000; B = 7'b1100010; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000000; B = 7'b1100010; | Outputs: P=%b | Expected: P=%d",
                 2329,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100111; B = 7'b0011001; // Expected: {'P': 2575}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100111; B = 7'b0011001; | Outputs: P=%b | Expected: P=%d",
                 2330,
                 
                 P
                 , 
                 
                 2575
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000101; B = 7'b1111110; // Expected: {'P': 8694}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000101; B = 7'b1111110; | Outputs: P=%b | Expected: P=%d",
                 2331,
                 
                 P
                 , 
                 
                 8694
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101110; B = 7'b1000111; // Expected: {'P': 7810}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101110; B = 7'b1000111; | Outputs: P=%b | Expected: P=%d",
                 2332,
                 
                 P
                 , 
                 
                 7810
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011101; B = 7'b1011000; // Expected: {'P': 2552}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011101; B = 7'b1011000; | Outputs: P=%b | Expected: P=%d",
                 2333,
                 
                 P
                 , 
                 
                 2552
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010100; B = 7'b1011000; // Expected: {'P': 1760}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010100; B = 7'b1011000; | Outputs: P=%b | Expected: P=%d",
                 2334,
                 
                 P
                 , 
                 
                 1760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001101; B = 7'b1011111; // Expected: {'P': 7315}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001101; B = 7'b1011111; | Outputs: P=%b | Expected: P=%d",
                 2335,
                 
                 P
                 , 
                 
                 7315
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100011; B = 7'b0010111; // Expected: {'P': 805}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100011; B = 7'b0010111; | Outputs: P=%b | Expected: P=%d",
                 2336,
                 
                 P
                 , 
                 
                 805
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000000; B = 7'b1001001; // Expected: {'P': 4672}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000000; B = 7'b1001001; | Outputs: P=%b | Expected: P=%d",
                 2337,
                 
                 P
                 , 
                 
                 4672
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001010; B = 7'b0010010; // Expected: {'P': 1332}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001010; B = 7'b0010010; | Outputs: P=%b | Expected: P=%d",
                 2338,
                 
                 P
                 , 
                 
                 1332
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011000; B = 7'b1110001; // Expected: {'P': 2712}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011000; B = 7'b1110001; | Outputs: P=%b | Expected: P=%d",
                 2339,
                 
                 P
                 , 
                 
                 2712
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001110; B = 7'b0100011; // Expected: {'P': 2730}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001110; B = 7'b0100011; | Outputs: P=%b | Expected: P=%d",
                 2340,
                 
                 P
                 , 
                 
                 2730
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101100; B = 7'b1000001; // Expected: {'P': 7020}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101100; B = 7'b1000001; | Outputs: P=%b | Expected: P=%d",
                 2341,
                 
                 P
                 , 
                 
                 7020
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111100; B = 7'b0011100; // Expected: {'P': 1680}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111100; B = 7'b0011100; | Outputs: P=%b | Expected: P=%d",
                 2342,
                 
                 P
                 , 
                 
                 1680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001000; B = 7'b1001000; // Expected: {'P': 576}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001000; B = 7'b1001000; | Outputs: P=%b | Expected: P=%d",
                 2343,
                 
                 P
                 , 
                 
                 576
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000010; B = 7'b1111001; // Expected: {'P': 7986}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000010; B = 7'b1111001; | Outputs: P=%b | Expected: P=%d",
                 2344,
                 
                 P
                 , 
                 
                 7986
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011010; B = 7'b0010011; // Expected: {'P': 1710}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011010; B = 7'b0010011; | Outputs: P=%b | Expected: P=%d",
                 2345,
                 
                 P
                 , 
                 
                 1710
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011001; B = 7'b0101000; // Expected: {'P': 3560}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011001; B = 7'b0101000; | Outputs: P=%b | Expected: P=%d",
                 2346,
                 
                 P
                 , 
                 
                 3560
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001011; B = 7'b1101001; // Expected: {'P': 7875}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001011; B = 7'b1101001; | Outputs: P=%b | Expected: P=%d",
                 2347,
                 
                 P
                 , 
                 
                 7875
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010011; B = 7'b1100010; // Expected: {'P': 8134}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010011; B = 7'b1100010; | Outputs: P=%b | Expected: P=%d",
                 2348,
                 
                 P
                 , 
                 
                 8134
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000101; B = 7'b0110101; // Expected: {'P': 265}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000101; B = 7'b0110101; | Outputs: P=%b | Expected: P=%d",
                 2349,
                 
                 P
                 , 
                 
                 265
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010010; B = 7'b1011110; // Expected: {'P': 7708}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010010; B = 7'b1011110; | Outputs: P=%b | Expected: P=%d",
                 2350,
                 
                 P
                 , 
                 
                 7708
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100011; B = 7'b0011111; // Expected: {'P': 1085}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100011; B = 7'b0011111; | Outputs: P=%b | Expected: P=%d",
                 2351,
                 
                 P
                 , 
                 
                 1085
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000000; B = 7'b1110001; // Expected: {'P': 7232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000000; B = 7'b1110001; | Outputs: P=%b | Expected: P=%d",
                 2352,
                 
                 P
                 , 
                 
                 7232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011000; B = 7'b0111101; // Expected: {'P': 1464}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011000; B = 7'b0111101; | Outputs: P=%b | Expected: P=%d",
                 2353,
                 
                 P
                 , 
                 
                 1464
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010101; B = 7'b0110110; // Expected: {'P': 1134}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010101; B = 7'b0110110; | Outputs: P=%b | Expected: P=%d",
                 2354,
                 
                 P
                 , 
                 
                 1134
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110100; B = 7'b0010000; // Expected: {'P': 832}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110100; B = 7'b0010000; | Outputs: P=%b | Expected: P=%d",
                 2355,
                 
                 P
                 , 
                 
                 832
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001011; B = 7'b0010011; // Expected: {'P': 209}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001011; B = 7'b0010011; | Outputs: P=%b | Expected: P=%d",
                 2356,
                 
                 P
                 , 
                 
                 209
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001101; B = 7'b1111011; // Expected: {'P': 9471}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001101; B = 7'b1111011; | Outputs: P=%b | Expected: P=%d",
                 2357,
                 
                 P
                 , 
                 
                 9471
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011100; B = 7'b1100111; // Expected: {'P': 9476}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011100; B = 7'b1100111; | Outputs: P=%b | Expected: P=%d",
                 2358,
                 
                 P
                 , 
                 
                 9476
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101011; B = 7'b0101011; // Expected: {'P': 4601}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101011; B = 7'b0101011; | Outputs: P=%b | Expected: P=%d",
                 2359,
                 
                 P
                 , 
                 
                 4601
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010101; B = 7'b0001000; // Expected: {'P': 680}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010101; B = 7'b0001000; | Outputs: P=%b | Expected: P=%d",
                 2360,
                 
                 P
                 , 
                 
                 680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001000; B = 7'b0011010; // Expected: {'P': 1872}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001000; B = 7'b0011010; | Outputs: P=%b | Expected: P=%d",
                 2361,
                 
                 P
                 , 
                 
                 1872
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100101; B = 7'b1011011; // Expected: {'P': 3367}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100101; B = 7'b1011011; | Outputs: P=%b | Expected: P=%d",
                 2362,
                 
                 P
                 , 
                 
                 3367
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100101; B = 7'b0110101; // Expected: {'P': 5353}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100101; B = 7'b0110101; | Outputs: P=%b | Expected: P=%d",
                 2363,
                 
                 P
                 , 
                 
                 5353
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010100; B = 7'b0100010; // Expected: {'P': 680}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010100; B = 7'b0100010; | Outputs: P=%b | Expected: P=%d",
                 2364,
                 
                 P
                 , 
                 
                 680
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111010; B = 7'b1100110; // Expected: {'P': 12444}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111010; B = 7'b1100110; | Outputs: P=%b | Expected: P=%d",
                 2365,
                 
                 P
                 , 
                 
                 12444
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111101; B = 7'b0001000; // Expected: {'P': 488}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111101; B = 7'b0001000; | Outputs: P=%b | Expected: P=%d",
                 2366,
                 
                 P
                 , 
                 
                 488
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010001; B = 7'b0100110; // Expected: {'P': 646}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010001; B = 7'b0100110; | Outputs: P=%b | Expected: P=%d",
                 2367,
                 
                 P
                 , 
                 
                 646
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110110; B = 7'b1010011; // Expected: {'P': 4482}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110110; B = 7'b1010011; | Outputs: P=%b | Expected: P=%d",
                 2368,
                 
                 P
                 , 
                 
                 4482
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011111; B = 7'b1011001; // Expected: {'P': 2759}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011111; B = 7'b1011001; | Outputs: P=%b | Expected: P=%d",
                 2369,
                 
                 P
                 , 
                 
                 2759
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110100; B = 7'b0000010; // Expected: {'P': 104}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110100; B = 7'b0000010; | Outputs: P=%b | Expected: P=%d",
                 2370,
                 
                 P
                 , 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001110; B = 7'b0010111; // Expected: {'P': 1794}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001110; B = 7'b0010111; | Outputs: P=%b | Expected: P=%d",
                 2371,
                 
                 P
                 , 
                 
                 1794
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111011; B = 7'b0110101; // Expected: {'P': 3127}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111011; B = 7'b0110101; | Outputs: P=%b | Expected: P=%d",
                 2372,
                 
                 P
                 , 
                 
                 3127
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110100; B = 7'b1010111; // Expected: {'P': 10092}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110100; B = 7'b1010111; | Outputs: P=%b | Expected: P=%d",
                 2373,
                 
                 P
                 , 
                 
                 10092
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010000; B = 7'b0101100; // Expected: {'P': 704}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010000; B = 7'b0101100; | Outputs: P=%b | Expected: P=%d",
                 2374,
                 
                 P
                 , 
                 
                 704
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011010; B = 7'b0001010; // Expected: {'P': 900}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011010; B = 7'b0001010; | Outputs: P=%b | Expected: P=%d",
                 2375,
                 
                 P
                 , 
                 
                 900
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110011; B = 7'b0010011; // Expected: {'P': 969}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110011; B = 7'b0010011; | Outputs: P=%b | Expected: P=%d",
                 2376,
                 
                 P
                 , 
                 
                 969
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111111; B = 7'b0111111; // Expected: {'P': 3969}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111111; B = 7'b0111111; | Outputs: P=%b | Expected: P=%d",
                 2377,
                 
                 P
                 , 
                 
                 3969
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001100; B = 7'b1111100; // Expected: {'P': 1488}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001100; B = 7'b1111100; | Outputs: P=%b | Expected: P=%d",
                 2378,
                 
                 P
                 , 
                 
                 1488
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001100; B = 7'b1110111; // Expected: {'P': 1428}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001100; B = 7'b1110111; | Outputs: P=%b | Expected: P=%d",
                 2379,
                 
                 P
                 , 
                 
                 1428
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101110; B = 7'b0010110; // Expected: {'P': 1012}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101110; B = 7'b0010110; | Outputs: P=%b | Expected: P=%d",
                 2380,
                 
                 P
                 , 
                 
                 1012
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111011; B = 7'b1011001; // Expected: {'P': 10947}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111011; B = 7'b1011001; | Outputs: P=%b | Expected: P=%d",
                 2381,
                 
                 P
                 , 
                 
                 10947
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100111; B = 7'b1010111; // Expected: {'P': 3393}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100111; B = 7'b1010111; | Outputs: P=%b | Expected: P=%d",
                 2382,
                 
                 P
                 , 
                 
                 3393
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111110; B = 7'b0011011; // Expected: {'P': 3402}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111110; B = 7'b0011011; | Outputs: P=%b | Expected: P=%d",
                 2383,
                 
                 P
                 , 
                 
                 3402
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110000; B = 7'b1111101; // Expected: {'P': 6000}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110000; B = 7'b1111101; | Outputs: P=%b | Expected: P=%d",
                 2384,
                 
                 P
                 , 
                 
                 6000
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010101; B = 7'b1010101; // Expected: {'P': 7225}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010101; B = 7'b1010101; | Outputs: P=%b | Expected: P=%d",
                 2385,
                 
                 P
                 , 
                 
                 7225
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100111; B = 7'b1000100; // Expected: {'P': 2652}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100111; B = 7'b1000100; | Outputs: P=%b | Expected: P=%d",
                 2386,
                 
                 P
                 , 
                 
                 2652
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110100; B = 7'b0011111; // Expected: {'P': 3596}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110100; B = 7'b0011111; | Outputs: P=%b | Expected: P=%d",
                 2387,
                 
                 P
                 , 
                 
                 3596
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000111; B = 7'b0001010; // Expected: {'P': 710}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000111; B = 7'b0001010; | Outputs: P=%b | Expected: P=%d",
                 2388,
                 
                 P
                 , 
                 
                 710
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110010; B = 7'b1000000; // Expected: {'P': 7296}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110010; B = 7'b1000000; | Outputs: P=%b | Expected: P=%d",
                 2389,
                 
                 P
                 , 
                 
                 7296
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010111; B = 7'b1101001; // Expected: {'P': 9135}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010111; B = 7'b1101001; | Outputs: P=%b | Expected: P=%d",
                 2390,
                 
                 P
                 , 
                 
                 9135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010001; B = 7'b1101011; // Expected: {'P': 8667}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010001; B = 7'b1101011; | Outputs: P=%b | Expected: P=%d",
                 2391,
                 
                 P
                 , 
                 
                 8667
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011110; B = 7'b0011011; // Expected: {'P': 810}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011110; B = 7'b0011011; | Outputs: P=%b | Expected: P=%d",
                 2392,
                 
                 P
                 , 
                 
                 810
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110110; B = 7'b0111001; // Expected: {'P': 3078}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110110; B = 7'b0111001; | Outputs: P=%b | Expected: P=%d",
                 2393,
                 
                 P
                 , 
                 
                 3078
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101000; B = 7'b0011100; // Expected: {'P': 1120}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101000; B = 7'b0011100; | Outputs: P=%b | Expected: P=%d",
                 2394,
                 
                 P
                 , 
                 
                 1120
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100010; B = 7'b0010101; // Expected: {'P': 2058}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100010; B = 7'b0010101; | Outputs: P=%b | Expected: P=%d",
                 2395,
                 
                 P
                 , 
                 
                 2058
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000111; B = 7'b1001000; // Expected: {'P': 504}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000111; B = 7'b1001000; | Outputs: P=%b | Expected: P=%d",
                 2396,
                 
                 P
                 , 
                 
                 504
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010111; B = 7'b1110001; // Expected: {'P': 9831}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010111; B = 7'b1110001; | Outputs: P=%b | Expected: P=%d",
                 2397,
                 
                 P
                 , 
                 
                 9831
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010100; B = 7'b0100111; // Expected: {'P': 780}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010100; B = 7'b0100111; | Outputs: P=%b | Expected: P=%d",
                 2398,
                 
                 P
                 , 
                 
                 780
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100000; B = 7'b0100001; // Expected: {'P': 3168}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100000; B = 7'b0100001; | Outputs: P=%b | Expected: P=%d",
                 2399,
                 
                 P
                 , 
                 
                 3168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010000; B = 7'b0010100; // Expected: {'P': 320}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010000; B = 7'b0010100; | Outputs: P=%b | Expected: P=%d",
                 2400,
                 
                 P
                 , 
                 
                 320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010001; B = 7'b1011011; // Expected: {'P': 1547}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010001; B = 7'b1011011; | Outputs: P=%b | Expected: P=%d",
                 2401,
                 
                 P
                 , 
                 
                 1547
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101101; B = 7'b0011110; // Expected: {'P': 1350}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101101; B = 7'b0011110; | Outputs: P=%b | Expected: P=%d",
                 2402,
                 
                 P
                 , 
                 
                 1350
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001100; B = 7'b0001110; // Expected: {'P': 168}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001100; B = 7'b0001110; | Outputs: P=%b | Expected: P=%d",
                 2403,
                 
                 P
                 , 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010001; B = 7'b0010101; // Expected: {'P': 1701}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010001; B = 7'b0010101; | Outputs: P=%b | Expected: P=%d",
                 2404,
                 
                 P
                 , 
                 
                 1701
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110011; B = 7'b1011000; // Expected: {'P': 4488}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110011; B = 7'b1011000; | Outputs: P=%b | Expected: P=%d",
                 2405,
                 
                 P
                 , 
                 
                 4488
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011010; B = 7'b0101001; // Expected: {'P': 1066}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011010; B = 7'b0101001; | Outputs: P=%b | Expected: P=%d",
                 2406,
                 
                 P
                 , 
                 
                 1066
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100111; B = 7'b1111111; // Expected: {'P': 13081}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100111; B = 7'b1111111; | Outputs: P=%b | Expected: P=%d",
                 2407,
                 
                 P
                 , 
                 
                 13081
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000000; B = 7'b0101100; // Expected: {'P': 2816}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000000; B = 7'b0101100; | Outputs: P=%b | Expected: P=%d",
                 2408,
                 
                 P
                 , 
                 
                 2816
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110111; B = 7'b0011001; // Expected: {'P': 2975}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110111; B = 7'b0011001; | Outputs: P=%b | Expected: P=%d",
                 2409,
                 
                 P
                 , 
                 
                 2975
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010001; B = 7'b1001010; // Expected: {'P': 5994}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010001; B = 7'b1001010; | Outputs: P=%b | Expected: P=%d",
                 2410,
                 
                 P
                 , 
                 
                 5994
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000000; B = 7'b1101100; // Expected: {'P': 6912}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000000; B = 7'b1101100; | Outputs: P=%b | Expected: P=%d",
                 2411,
                 
                 P
                 , 
                 
                 6912
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001110; B = 7'b0101111; // Expected: {'P': 3666}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001110; B = 7'b0101111; | Outputs: P=%b | Expected: P=%d",
                 2412,
                 
                 P
                 , 
                 
                 3666
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101100; B = 7'b0001000; // Expected: {'P': 352}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101100; B = 7'b0001000; | Outputs: P=%b | Expected: P=%d",
                 2413,
                 
                 P
                 , 
                 
                 352
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110111; B = 7'b1100101; // Expected: {'P': 5555}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110111; B = 7'b1100101; | Outputs: P=%b | Expected: P=%d",
                 2414,
                 
                 P
                 , 
                 
                 5555
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000000; B = 7'b1011111; // Expected: {'P': 6080}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000000; B = 7'b1011111; | Outputs: P=%b | Expected: P=%d",
                 2415,
                 
                 P
                 , 
                 
                 6080
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110111; B = 7'b1011101; // Expected: {'P': 11067}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110111; B = 7'b1011101; | Outputs: P=%b | Expected: P=%d",
                 2416,
                 
                 P
                 , 
                 
                 11067
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010100; B = 7'b1011010; // Expected: {'P': 1800}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010100; B = 7'b1011010; | Outputs: P=%b | Expected: P=%d",
                 2417,
                 
                 P
                 , 
                 
                 1800
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111110; B = 7'b1010100; // Expected: {'P': 5208}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111110; B = 7'b1010100; | Outputs: P=%b | Expected: P=%d",
                 2418,
                 
                 P
                 , 
                 
                 5208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011000; B = 7'b0100000; // Expected: {'P': 2816}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011000; B = 7'b0100000; | Outputs: P=%b | Expected: P=%d",
                 2419,
                 
                 P
                 , 
                 
                 2816
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001100; B = 7'b0100001; // Expected: {'P': 2508}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001100; B = 7'b0100001; | Outputs: P=%b | Expected: P=%d",
                 2420,
                 
                 P
                 , 
                 
                 2508
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000011; B = 7'b1101000; // Expected: {'P': 312}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000011; B = 7'b1101000; | Outputs: P=%b | Expected: P=%d",
                 2421,
                 
                 P
                 , 
                 
                 312
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110011; B = 7'b0101100; // Expected: {'P': 5060}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110011; B = 7'b0101100; | Outputs: P=%b | Expected: P=%d",
                 2422,
                 
                 P
                 , 
                 
                 5060
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101100; B = 7'b0110010; // Expected: {'P': 2200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101100; B = 7'b0110010; | Outputs: P=%b | Expected: P=%d",
                 2423,
                 
                 P
                 , 
                 
                 2200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100010; B = 7'b1000010; // Expected: {'P': 2244}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100010; B = 7'b1000010; | Outputs: P=%b | Expected: P=%d",
                 2424,
                 
                 P
                 , 
                 
                 2244
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011100; B = 7'b0000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011100; B = 7'b0000000; | Outputs: P=%b | Expected: P=%d",
                 2425,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011011; B = 7'b1111111; // Expected: {'P': 11557}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011011; B = 7'b1111111; | Outputs: P=%b | Expected: P=%d",
                 2426,
                 
                 P
                 , 
                 
                 11557
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100010; B = 7'b1110010; // Expected: {'P': 3876}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100010; B = 7'b1110010; | Outputs: P=%b | Expected: P=%d",
                 2427,
                 
                 P
                 , 
                 
                 3876
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010101; B = 7'b1011100; // Expected: {'P': 7820}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010101; B = 7'b1011100; | Outputs: P=%b | Expected: P=%d",
                 2428,
                 
                 P
                 , 
                 
                 7820
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011110; B = 7'b1111001; // Expected: {'P': 3630}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011110; B = 7'b1111001; | Outputs: P=%b | Expected: P=%d",
                 2429,
                 
                 P
                 , 
                 
                 3630
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001110; B = 7'b1000101; // Expected: {'P': 966}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001110; B = 7'b1000101; | Outputs: P=%b | Expected: P=%d",
                 2430,
                 
                 P
                 , 
                 
                 966
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001100; B = 7'b0110101; // Expected: {'P': 4028}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001100; B = 7'b0110101; | Outputs: P=%b | Expected: P=%d",
                 2431,
                 
                 P
                 , 
                 
                 4028
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100111; B = 7'b1001111; // Expected: {'P': 8137}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100111; B = 7'b1001111; | Outputs: P=%b | Expected: P=%d",
                 2432,
                 
                 P
                 , 
                 
                 8137
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100110; B = 7'b0101111; // Expected: {'P': 1786}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100110; B = 7'b0101111; | Outputs: P=%b | Expected: P=%d",
                 2433,
                 
                 P
                 , 
                 
                 1786
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000010; B = 7'b1010000; // Expected: {'P': 160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000010; B = 7'b1010000; | Outputs: P=%b | Expected: P=%d",
                 2434,
                 
                 P
                 , 
                 
                 160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001110; B = 7'b1101001; // Expected: {'P': 8190}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001110; B = 7'b1101001; | Outputs: P=%b | Expected: P=%d",
                 2435,
                 
                 P
                 , 
                 
                 8190
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000101; B = 7'b1001111; // Expected: {'P': 5451}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000101; B = 7'b1001111; | Outputs: P=%b | Expected: P=%d",
                 2436,
                 
                 P
                 , 
                 
                 5451
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111110; B = 7'b0101110; // Expected: {'P': 2852}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111110; B = 7'b0101110; | Outputs: P=%b | Expected: P=%d",
                 2437,
                 
                 P
                 , 
                 
                 2852
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100101; B = 7'b0010000; // Expected: {'P': 1616}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100101; B = 7'b0010000; | Outputs: P=%b | Expected: P=%d",
                 2438,
                 
                 P
                 , 
                 
                 1616
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011101; B = 7'b0101000; // Expected: {'P': 1160}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011101; B = 7'b0101000; | Outputs: P=%b | Expected: P=%d",
                 2439,
                 
                 P
                 , 
                 
                 1160
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111111; B = 7'b1010010; // Expected: {'P': 10414}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111111; B = 7'b1010010; | Outputs: P=%b | Expected: P=%d",
                 2440,
                 
                 P
                 , 
                 
                 10414
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101100; B = 7'b0000001; // Expected: {'P': 108}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101100; B = 7'b0000001; | Outputs: P=%b | Expected: P=%d",
                 2441,
                 
                 P
                 , 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011011; B = 7'b1001001; // Expected: {'P': 6643}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011011; B = 7'b1001001; | Outputs: P=%b | Expected: P=%d",
                 2442,
                 
                 P
                 , 
                 
                 6643
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101100; B = 7'b1001000; // Expected: {'P': 3168}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101100; B = 7'b1001000; | Outputs: P=%b | Expected: P=%d",
                 2443,
                 
                 P
                 , 
                 
                 3168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010000; B = 7'b0000001; // Expected: {'P': 80}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010000; B = 7'b0000001; | Outputs: P=%b | Expected: P=%d",
                 2444,
                 
                 P
                 , 
                 
                 80
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000000; B = 7'b0110010; // Expected: {'P': 3200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000000; B = 7'b0110010; | Outputs: P=%b | Expected: P=%d",
                 2445,
                 
                 P
                 , 
                 
                 3200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000000; B = 7'b0001101; // Expected: {'P': 832}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000000; B = 7'b0001101; | Outputs: P=%b | Expected: P=%d",
                 2446,
                 
                 P
                 , 
                 
                 832
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001011; B = 7'b1110100; // Expected: {'P': 8700}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001011; B = 7'b1110100; | Outputs: P=%b | Expected: P=%d",
                 2447,
                 
                 P
                 , 
                 
                 8700
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000101; B = 7'b1011010; // Expected: {'P': 450}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000101; B = 7'b1011010; | Outputs: P=%b | Expected: P=%d",
                 2448,
                 
                 P
                 , 
                 
                 450
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001101; B = 7'b1101011; // Expected: {'P': 8239}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001101; B = 7'b1101011; | Outputs: P=%b | Expected: P=%d",
                 2449,
                 
                 P
                 , 
                 
                 8239
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010100; B = 7'b1000001; // Expected: {'P': 1300}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010100; B = 7'b1000001; | Outputs: P=%b | Expected: P=%d",
                 2450,
                 
                 P
                 , 
                 
                 1300
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010111; B = 7'b0100000; // Expected: {'P': 736}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010111; B = 7'b0100000; | Outputs: P=%b | Expected: P=%d",
                 2451,
                 
                 P
                 , 
                 
                 736
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101101; B = 7'b0000110; // Expected: {'P': 654}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101101; B = 7'b0000110; | Outputs: P=%b | Expected: P=%d",
                 2452,
                 
                 P
                 , 
                 
                 654
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101100; B = 7'b1000011; // Expected: {'P': 7236}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101100; B = 7'b1000011; | Outputs: P=%b | Expected: P=%d",
                 2453,
                 
                 P
                 , 
                 
                 7236
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111010; B = 7'b1001001; // Expected: {'P': 4234}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111010; B = 7'b1001001; | Outputs: P=%b | Expected: P=%d",
                 2454,
                 
                 P
                 , 
                 
                 4234
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101010; B = 7'b1000011; // Expected: {'P': 2814}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101010; B = 7'b1000011; | Outputs: P=%b | Expected: P=%d",
                 2455,
                 
                 P
                 , 
                 
                 2814
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011101; B = 7'b1101000; // Expected: {'P': 9672}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011101; B = 7'b1101000; | Outputs: P=%b | Expected: P=%d",
                 2456,
                 
                 P
                 , 
                 
                 9672
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000111; B = 7'b0110101; // Expected: {'P': 371}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000111; B = 7'b0110101; | Outputs: P=%b | Expected: P=%d",
                 2457,
                 
                 P
                 , 
                 
                 371
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111100; B = 7'b1110111; // Expected: {'P': 14756}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111100; B = 7'b1110111; | Outputs: P=%b | Expected: P=%d",
                 2458,
                 
                 P
                 , 
                 
                 14756
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010101; B = 7'b0010111; // Expected: {'P': 1955}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010101; B = 7'b0010111; | Outputs: P=%b | Expected: P=%d",
                 2459,
                 
                 P
                 , 
                 
                 1955
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111000; B = 7'b1011010; // Expected: {'P': 5040}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111000; B = 7'b1011010; | Outputs: P=%b | Expected: P=%d",
                 2460,
                 
                 P
                 , 
                 
                 5040
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110110; B = 7'b0000011; // Expected: {'P': 162}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110110; B = 7'b0000011; | Outputs: P=%b | Expected: P=%d",
                 2461,
                 
                 P
                 , 
                 
                 162
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001011; B = 7'b1000110; // Expected: {'P': 770}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001011; B = 7'b1000110; | Outputs: P=%b | Expected: P=%d",
                 2462,
                 
                 P
                 , 
                 
                 770
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000001; B = 7'b1110110; // Expected: {'P': 7670}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000001; B = 7'b1110110; | Outputs: P=%b | Expected: P=%d",
                 2463,
                 
                 P
                 , 
                 
                 7670
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110001; B = 7'b0001101; // Expected: {'P': 1469}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110001; B = 7'b0001101; | Outputs: P=%b | Expected: P=%d",
                 2464,
                 
                 P
                 , 
                 
                 1469
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101010; B = 7'b1101111; // Expected: {'P': 11766}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101010; B = 7'b1101111; | Outputs: P=%b | Expected: P=%d",
                 2465,
                 
                 P
                 , 
                 
                 11766
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110111; B = 7'b1001000; // Expected: {'P': 3960}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110111; B = 7'b1001000; | Outputs: P=%b | Expected: P=%d",
                 2466,
                 
                 P
                 , 
                 
                 3960
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101010; B = 7'b1011101; // Expected: {'P': 9858}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101010; B = 7'b1011101; | Outputs: P=%b | Expected: P=%d",
                 2467,
                 
                 P
                 , 
                 
                 9858
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010001; B = 7'b0001110; // Expected: {'P': 1134}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010001; B = 7'b0001110; | Outputs: P=%b | Expected: P=%d",
                 2468,
                 
                 P
                 , 
                 
                 1134
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000001; B = 7'b1101000; // Expected: {'P': 104}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000001; B = 7'b1101000; | Outputs: P=%b | Expected: P=%d",
                 2469,
                 
                 P
                 , 
                 
                 104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001110; B = 7'b1001001; // Expected: {'P': 5694}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001110; B = 7'b1001001; | Outputs: P=%b | Expected: P=%d",
                 2470,
                 
                 P
                 , 
                 
                 5694
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100111; B = 7'b0001001; // Expected: {'P': 351}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100111; B = 7'b0001001; | Outputs: P=%b | Expected: P=%d",
                 2471,
                 
                 P
                 , 
                 
                 351
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101110; B = 7'b0111011; // Expected: {'P': 6490}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101110; B = 7'b0111011; | Outputs: P=%b | Expected: P=%d",
                 2472,
                 
                 P
                 , 
                 
                 6490
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010011; B = 7'b1001000; // Expected: {'P': 5976}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010011; B = 7'b1001000; | Outputs: P=%b | Expected: P=%d",
                 2473,
                 
                 P
                 , 
                 
                 5976
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000001; B = 7'b0001111; // Expected: {'P': 975}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000001; B = 7'b0001111; | Outputs: P=%b | Expected: P=%d",
                 2474,
                 
                 P
                 , 
                 
                 975
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111100; B = 7'b0111110; // Expected: {'P': 7688}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111100; B = 7'b0111110; | Outputs: P=%b | Expected: P=%d",
                 2475,
                 
                 P
                 , 
                 
                 7688
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111001; B = 7'b1011000; // Expected: {'P': 10648}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111001; B = 7'b1011000; | Outputs: P=%b | Expected: P=%d",
                 2476,
                 
                 P
                 , 
                 
                 10648
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110110; B = 7'b0010010; // Expected: {'P': 2124}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110110; B = 7'b0010010; | Outputs: P=%b | Expected: P=%d",
                 2477,
                 
                 P
                 , 
                 
                 2124
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000010; B = 7'b0101111; // Expected: {'P': 94}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000010; B = 7'b0101111; | Outputs: P=%b | Expected: P=%d",
                 2478,
                 
                 P
                 , 
                 
                 94
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111110; B = 7'b1110001; // Expected: {'P': 14238}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111110; B = 7'b1110001; | Outputs: P=%b | Expected: P=%d",
                 2479,
                 
                 P
                 , 
                 
                 14238
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111101; B = 7'b1011001; // Expected: {'P': 11125}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111101; B = 7'b1011001; | Outputs: P=%b | Expected: P=%d",
                 2480,
                 
                 P
                 , 
                 
                 11125
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111111; B = 7'b0001000; // Expected: {'P': 1016}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111111; B = 7'b0001000; | Outputs: P=%b | Expected: P=%d",
                 2481,
                 
                 P
                 , 
                 
                 1016
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011000; B = 7'b0111111; // Expected: {'P': 1512}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011000; B = 7'b0111111; | Outputs: P=%b | Expected: P=%d",
                 2482,
                 
                 P
                 , 
                 
                 1512
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011000; B = 7'b1110000; // Expected: {'P': 9856}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011000; B = 7'b1110000; | Outputs: P=%b | Expected: P=%d",
                 2483,
                 
                 P
                 , 
                 
                 9856
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000000; B = 7'b1001111; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000000; B = 7'b1001111; | Outputs: P=%b | Expected: P=%d",
                 2484,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001011; B = 7'b1001010; // Expected: {'P': 5550}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001011; B = 7'b1001010; | Outputs: P=%b | Expected: P=%d",
                 2485,
                 
                 P
                 , 
                 
                 5550
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011111; B = 7'b0111101; // Expected: {'P': 1891}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011111; B = 7'b0111101; | Outputs: P=%b | Expected: P=%d",
                 2486,
                 
                 P
                 , 
                 
                 1891
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100101; B = 7'b0011111; // Expected: {'P': 3131}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100101; B = 7'b0011111; | Outputs: P=%b | Expected: P=%d",
                 2487,
                 
                 P
                 , 
                 
                 3131
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100011; B = 7'b0111110; // Expected: {'P': 6138}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100011; B = 7'b0111110; | Outputs: P=%b | Expected: P=%d",
                 2488,
                 
                 P
                 , 
                 
                 6138
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100011; B = 7'b1010000; // Expected: {'P': 7920}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100011; B = 7'b1010000; | Outputs: P=%b | Expected: P=%d",
                 2489,
                 
                 P
                 , 
                 
                 7920
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010001; B = 7'b1101100; // Expected: {'P': 8748}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010001; B = 7'b1101100; | Outputs: P=%b | Expected: P=%d",
                 2490,
                 
                 P
                 , 
                 
                 8748
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101110; B = 7'b1101000; // Expected: {'P': 4784}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101110; B = 7'b1101000; | Outputs: P=%b | Expected: P=%d",
                 2491,
                 
                 P
                 , 
                 
                 4784
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110100; B = 7'b1111010; // Expected: {'P': 6344}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110100; B = 7'b1111010; | Outputs: P=%b | Expected: P=%d",
                 2492,
                 
                 P
                 , 
                 
                 6344
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100011; B = 7'b1111010; // Expected: {'P': 12078}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100011; B = 7'b1111010; | Outputs: P=%b | Expected: P=%d",
                 2493,
                 
                 P
                 , 
                 
                 12078
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001000; B = 7'b1101111; // Expected: {'P': 888}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001000; B = 7'b1101111; | Outputs: P=%b | Expected: P=%d",
                 2494,
                 
                 P
                 , 
                 
                 888
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101110; B = 7'b1000001; // Expected: {'P': 2990}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101110; B = 7'b1000001; | Outputs: P=%b | Expected: P=%d",
                 2495,
                 
                 P
                 , 
                 
                 2990
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010001; B = 7'b1011001; // Expected: {'P': 7209}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010001; B = 7'b1011001; | Outputs: P=%b | Expected: P=%d",
                 2496,
                 
                 P
                 , 
                 
                 7209
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010111; B = 7'b1011011; // Expected: {'P': 2093}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010111; B = 7'b1011011; | Outputs: P=%b | Expected: P=%d",
                 2497,
                 
                 P
                 , 
                 
                 2093
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010101; B = 7'b1010010; // Expected: {'P': 6970}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010101; B = 7'b1010010; | Outputs: P=%b | Expected: P=%d",
                 2498,
                 
                 P
                 , 
                 
                 6970
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100111; B = 7'b1010110; // Expected: {'P': 8858}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100111; B = 7'b1010110; | Outputs: P=%b | Expected: P=%d",
                 2499,
                 
                 P
                 , 
                 
                 8858
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100101; B = 7'b1101101; // Expected: {'P': 11009}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100101; B = 7'b1101101; | Outputs: P=%b | Expected: P=%d",
                 2500,
                 
                 P
                 , 
                 
                 11009
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111001; B = 7'b1101110; // Expected: {'P': 13310}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111001; B = 7'b1101110; | Outputs: P=%b | Expected: P=%d",
                 2501,
                 
                 P
                 , 
                 
                 13310
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101111; B = 7'b0111001; // Expected: {'P': 6327}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101111; B = 7'b0111001; | Outputs: P=%b | Expected: P=%d",
                 2502,
                 
                 P
                 , 
                 
                 6327
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101111; B = 7'b0010110; // Expected: {'P': 2442}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101111; B = 7'b0010110; | Outputs: P=%b | Expected: P=%d",
                 2503,
                 
                 P
                 , 
                 
                 2442
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110111; B = 7'b0011110; // Expected: {'P': 1650}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110111; B = 7'b0011110; | Outputs: P=%b | Expected: P=%d",
                 2504,
                 
                 P
                 , 
                 
                 1650
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111010; B = 7'b1100010; // Expected: {'P': 5684}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111010; B = 7'b1100010; | Outputs: P=%b | Expected: P=%d",
                 2505,
                 
                 P
                 , 
                 
                 5684
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010111; B = 7'b0111010; // Expected: {'P': 1334}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010111; B = 7'b0111010; | Outputs: P=%b | Expected: P=%d",
                 2506,
                 
                 P
                 , 
                 
                 1334
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100011; B = 7'b1111111; // Expected: {'P': 12573}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100011; B = 7'b1111111; | Outputs: P=%b | Expected: P=%d",
                 2507,
                 
                 P
                 , 
                 
                 12573
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100001; B = 7'b0010101; // Expected: {'P': 2037}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100001; B = 7'b0010101; | Outputs: P=%b | Expected: P=%d",
                 2508,
                 
                 P
                 , 
                 
                 2037
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111101; B = 7'b1100111; // Expected: {'P': 12875}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111101; B = 7'b1100111; | Outputs: P=%b | Expected: P=%d",
                 2509,
                 
                 P
                 , 
                 
                 12875
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000111; B = 7'b1001001; // Expected: {'P': 5183}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000111; B = 7'b1001001; | Outputs: P=%b | Expected: P=%d",
                 2510,
                 
                 P
                 , 
                 
                 5183
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101011; B = 7'b1101011; // Expected: {'P': 4601}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101011; B = 7'b1101011; | Outputs: P=%b | Expected: P=%d",
                 2511,
                 
                 P
                 , 
                 
                 4601
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000000; B = 7'b1010111; // Expected: {'P': 5568}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000000; B = 7'b1010111; | Outputs: P=%b | Expected: P=%d",
                 2512,
                 
                 P
                 , 
                 
                 5568
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000010; B = 7'b0011101; // Expected: {'P': 1914}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000010; B = 7'b0011101; | Outputs: P=%b | Expected: P=%d",
                 2513,
                 
                 P
                 , 
                 
                 1914
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101010; B = 7'b0010111; // Expected: {'P': 966}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101010; B = 7'b0010111; | Outputs: P=%b | Expected: P=%d",
                 2514,
                 
                 P
                 , 
                 
                 966
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001000; B = 7'b0011101; // Expected: {'P': 2088}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001000; B = 7'b0011101; | Outputs: P=%b | Expected: P=%d",
                 2515,
                 
                 P
                 , 
                 
                 2088
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111011; B = 7'b0001010; // Expected: {'P': 590}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111011; B = 7'b0001010; | Outputs: P=%b | Expected: P=%d",
                 2516,
                 
                 P
                 , 
                 
                 590
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101010; B = 7'b0111101; // Expected: {'P': 2562}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101010; B = 7'b0111101; | Outputs: P=%b | Expected: P=%d",
                 2517,
                 
                 P
                 , 
                 
                 2562
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100100; B = 7'b1011000; // Expected: {'P': 3168}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100100; B = 7'b1011000; | Outputs: P=%b | Expected: P=%d",
                 2518,
                 
                 P
                 , 
                 
                 3168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010100; B = 7'b1010110; // Expected: {'P': 1720}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010100; B = 7'b1010110; | Outputs: P=%b | Expected: P=%d",
                 2519,
                 
                 P
                 , 
                 
                 1720
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001110; B = 7'b0010001; // Expected: {'P': 1326}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001110; B = 7'b0010001; | Outputs: P=%b | Expected: P=%d",
                 2520,
                 
                 P
                 , 
                 
                 1326
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100100; B = 7'b0111000; // Expected: {'P': 5600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100100; B = 7'b0111000; | Outputs: P=%b | Expected: P=%d",
                 2521,
                 
                 P
                 , 
                 
                 5600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001110; B = 7'b0111001; // Expected: {'P': 4446}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001110; B = 7'b0111001; | Outputs: P=%b | Expected: P=%d",
                 2522,
                 
                 P
                 , 
                 
                 4446
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000101; B = 7'b1010000; // Expected: {'P': 400}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000101; B = 7'b1010000; | Outputs: P=%b | Expected: P=%d",
                 2523,
                 
                 P
                 , 
                 
                 400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100101; B = 7'b0111001; // Expected: {'P': 5757}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100101; B = 7'b0111001; | Outputs: P=%b | Expected: P=%d",
                 2524,
                 
                 P
                 , 
                 
                 5757
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100000; B = 7'b0111100; // Expected: {'P': 5760}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100000; B = 7'b0111100; | Outputs: P=%b | Expected: P=%d",
                 2525,
                 
                 P
                 , 
                 
                 5760
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101111; B = 7'b1111010; // Expected: {'P': 13542}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101111; B = 7'b1111010; | Outputs: P=%b | Expected: P=%d",
                 2526,
                 
                 P
                 , 
                 
                 13542
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011011; B = 7'b1010111; // Expected: {'P': 2349}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011011; B = 7'b1010111; | Outputs: P=%b | Expected: P=%d",
                 2527,
                 
                 P
                 , 
                 
                 2349
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011101; B = 7'b1000011; // Expected: {'P': 1943}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011101; B = 7'b1000011; | Outputs: P=%b | Expected: P=%d",
                 2528,
                 
                 P
                 , 
                 
                 1943
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000000; B = 7'b1100001; // Expected: {'P': 6208}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000000; B = 7'b1100001; | Outputs: P=%b | Expected: P=%d",
                 2529,
                 
                 P
                 , 
                 
                 6208
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110101; B = 7'b1111111; // Expected: {'P': 14859}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110101; B = 7'b1111111; | Outputs: P=%b | Expected: P=%d",
                 2530,
                 
                 P
                 , 
                 
                 14859
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111110; B = 7'b1001000; // Expected: {'P': 4464}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111110; B = 7'b1001000; | Outputs: P=%b | Expected: P=%d",
                 2531,
                 
                 P
                 , 
                 
                 4464
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101001; B = 7'b1100001; // Expected: {'P': 3977}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101001; B = 7'b1100001; | Outputs: P=%b | Expected: P=%d",
                 2532,
                 
                 P
                 , 
                 
                 3977
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001010; B = 7'b0110110; // Expected: {'P': 3996}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001010; B = 7'b0110110; | Outputs: P=%b | Expected: P=%d",
                 2533,
                 
                 P
                 , 
                 
                 3996
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111100; B = 7'b0110011; // Expected: {'P': 3060}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111100; B = 7'b0110011; | Outputs: P=%b | Expected: P=%d",
                 2534,
                 
                 P
                 , 
                 
                 3060
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100001; B = 7'b0100000; // Expected: {'P': 3104}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100001; B = 7'b0100000; | Outputs: P=%b | Expected: P=%d",
                 2535,
                 
                 P
                 , 
                 
                 3104
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101100; B = 7'b1001110; // Expected: {'P': 8424}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101100; B = 7'b1001110; | Outputs: P=%b | Expected: P=%d",
                 2536,
                 
                 P
                 , 
                 
                 8424
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011000; B = 7'b1010110; // Expected: {'P': 7568}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011000; B = 7'b1010110; | Outputs: P=%b | Expected: P=%d",
                 2537,
                 
                 P
                 , 
                 
                 7568
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010101; B = 7'b0001011; // Expected: {'P': 231}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010101; B = 7'b0001011; | Outputs: P=%b | Expected: P=%d",
                 2538,
                 
                 P
                 , 
                 
                 231
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111111; B = 7'b1011001; // Expected: {'P': 11303}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111111; B = 7'b1011001; | Outputs: P=%b | Expected: P=%d",
                 2539,
                 
                 P
                 , 
                 
                 11303
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000010; B = 7'b1000011; // Expected: {'P': 134}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000010; B = 7'b1000011; | Outputs: P=%b | Expected: P=%d",
                 2540,
                 
                 P
                 , 
                 
                 134
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111101; B = 7'b0000111; // Expected: {'P': 875}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111101; B = 7'b0000111; | Outputs: P=%b | Expected: P=%d",
                 2541,
                 
                 P
                 , 
                 
                 875
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101100; B = 7'b0111011; // Expected: {'P': 2596}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101100; B = 7'b0111011; | Outputs: P=%b | Expected: P=%d",
                 2542,
                 
                 P
                 , 
                 
                 2596
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110011; B = 7'b0001111; // Expected: {'P': 765}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110011; B = 7'b0001111; | Outputs: P=%b | Expected: P=%d",
                 2543,
                 
                 P
                 , 
                 
                 765
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110111; B = 7'b1000010; // Expected: {'P': 3630}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110111; B = 7'b1000010; | Outputs: P=%b | Expected: P=%d",
                 2544,
                 
                 P
                 , 
                 
                 3630
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111110; B = 7'b0101000; // Expected: {'P': 2480}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111110; B = 7'b0101000; | Outputs: P=%b | Expected: P=%d",
                 2545,
                 
                 P
                 , 
                 
                 2480
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110110; B = 7'b1100000; // Expected: {'P': 5184}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110110; B = 7'b1100000; | Outputs: P=%b | Expected: P=%d",
                 2546,
                 
                 P
                 , 
                 
                 5184
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000010; B = 7'b0011001; // Expected: {'P': 1650}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000010; B = 7'b0011001; | Outputs: P=%b | Expected: P=%d",
                 2547,
                 
                 P
                 , 
                 
                 1650
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101111; B = 7'b1100011; // Expected: {'P': 10989}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101111; B = 7'b1100011; | Outputs: P=%b | Expected: P=%d",
                 2548,
                 
                 P
                 , 
                 
                 10989
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010010; B = 7'b0100010; // Expected: {'P': 2788}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010010; B = 7'b0100010; | Outputs: P=%b | Expected: P=%d",
                 2549,
                 
                 P
                 , 
                 
                 2788
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101110; B = 7'b0110111; // Expected: {'P': 6050}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101110; B = 7'b0110111; | Outputs: P=%b | Expected: P=%d",
                 2550,
                 
                 P
                 , 
                 
                 6050
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000110; B = 7'b1000000; // Expected: {'P': 384}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000110; B = 7'b1000000; | Outputs: P=%b | Expected: P=%d",
                 2551,
                 
                 P
                 , 
                 
                 384
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011111; B = 7'b1110101; // Expected: {'P': 3627}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011111; B = 7'b1110101; | Outputs: P=%b | Expected: P=%d",
                 2552,
                 
                 P
                 , 
                 
                 3627
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101101; B = 7'b1101100; // Expected: {'P': 4860}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101101; B = 7'b1101100; | Outputs: P=%b | Expected: P=%d",
                 2553,
                 
                 P
                 , 
                 
                 4860
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111001; B = 7'b0010011; // Expected: {'P': 1083}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111001; B = 7'b0010011; | Outputs: P=%b | Expected: P=%d",
                 2554,
                 
                 P
                 , 
                 
                 1083
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101111; B = 7'b0101100; // Expected: {'P': 4884}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101111; B = 7'b0101100; | Outputs: P=%b | Expected: P=%d",
                 2555,
                 
                 P
                 , 
                 
                 4884
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111010; B = 7'b0001101; // Expected: {'P': 1586}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111010; B = 7'b0001101; | Outputs: P=%b | Expected: P=%d",
                 2556,
                 
                 P
                 , 
                 
                 1586
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101000; B = 7'b0100001; // Expected: {'P': 1320}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101000; B = 7'b0100001; | Outputs: P=%b | Expected: P=%d",
                 2557,
                 
                 P
                 , 
                 
                 1320
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000001; B = 7'b0111000; // Expected: {'P': 56}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000001; B = 7'b0111000; | Outputs: P=%b | Expected: P=%d",
                 2558,
                 
                 P
                 , 
                 
                 56
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011000; B = 7'b1100111; // Expected: {'P': 2472}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011000; B = 7'b1100111; | Outputs: P=%b | Expected: P=%d",
                 2559,
                 
                 P
                 , 
                 
                 2472
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011000; B = 7'b0010111; // Expected: {'P': 2024}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011000; B = 7'b0010111; | Outputs: P=%b | Expected: P=%d",
                 2560,
                 
                 P
                 , 
                 
                 2024
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000111; B = 7'b0000001; // Expected: {'P': 7}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000111; B = 7'b0000001; | Outputs: P=%b | Expected: P=%d",
                 2561,
                 
                 P
                 , 
                 
                 7
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101000; B = 7'b0001110; // Expected: {'P': 1456}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101000; B = 7'b0001110; | Outputs: P=%b | Expected: P=%d",
                 2562,
                 
                 P
                 , 
                 
                 1456
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010000; B = 7'b0000000; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010000; B = 7'b0000000; | Outputs: P=%b | Expected: P=%d",
                 2563,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100101; B = 7'b0101101; // Expected: {'P': 4545}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100101; B = 7'b0101101; | Outputs: P=%b | Expected: P=%d",
                 2564,
                 
                 P
                 , 
                 
                 4545
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100111; B = 7'b0001110; // Expected: {'P': 546}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100111; B = 7'b0001110; | Outputs: P=%b | Expected: P=%d",
                 2565,
                 
                 P
                 , 
                 
                 546
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110111; B = 7'b1111010; // Expected: {'P': 6710}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110111; B = 7'b1111010; | Outputs: P=%b | Expected: P=%d",
                 2566,
                 
                 P
                 , 
                 
                 6710
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100101; B = 7'b0001000; // Expected: {'P': 808}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100101; B = 7'b0001000; | Outputs: P=%b | Expected: P=%d",
                 2567,
                 
                 P
                 , 
                 
                 808
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000101; B = 7'b0000111; // Expected: {'P': 483}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000101; B = 7'b0000111; | Outputs: P=%b | Expected: P=%d",
                 2568,
                 
                 P
                 , 
                 
                 483
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100111; B = 7'b1100110; // Expected: {'P': 10506}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100111; B = 7'b1100110; | Outputs: P=%b | Expected: P=%d",
                 2569,
                 
                 P
                 , 
                 
                 10506
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010000; B = 7'b0010110; // Expected: {'P': 352}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010000; B = 7'b0010110; | Outputs: P=%b | Expected: P=%d",
                 2570,
                 
                 P
                 , 
                 
                 352
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011110; B = 7'b0101111; // Expected: {'P': 4418}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011110; B = 7'b0101111; | Outputs: P=%b | Expected: P=%d",
                 2571,
                 
                 P
                 , 
                 
                 4418
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1101010; B = 7'b0001000; // Expected: {'P': 848}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1101010; B = 7'b0001000; | Outputs: P=%b | Expected: P=%d",
                 2572,
                 
                 P
                 , 
                 
                 848
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000101; B = 7'b1000000; // Expected: {'P': 4416}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000101; B = 7'b1000000; | Outputs: P=%b | Expected: P=%d",
                 2573,
                 
                 P
                 , 
                 
                 4416
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011000; B = 7'b1001111; // Expected: {'P': 6952}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011000; B = 7'b1001111; | Outputs: P=%b | Expected: P=%d",
                 2574,
                 
                 P
                 , 
                 
                 6952
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001000; B = 7'b0011101; // Expected: {'P': 232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001000; B = 7'b0011101; | Outputs: P=%b | Expected: P=%d",
                 2575,
                 
                 P
                 , 
                 
                 232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000011; B = 7'b0100100; // Expected: {'P': 108}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000011; B = 7'b0100100; | Outputs: P=%b | Expected: P=%d",
                 2576,
                 
                 P
                 , 
                 
                 108
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000010; B = 7'b1110101; // Expected: {'P': 234}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000010; B = 7'b1110101; | Outputs: P=%b | Expected: P=%d",
                 2577,
                 
                 P
                 , 
                 
                 234
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011000; B = 7'b0001100; // Expected: {'P': 288}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011000; B = 7'b0001100; | Outputs: P=%b | Expected: P=%d",
                 2578,
                 
                 P
                 , 
                 
                 288
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100010; B = 7'b0101111; // Expected: {'P': 4606}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100010; B = 7'b0101111; | Outputs: P=%b | Expected: P=%d",
                 2579,
                 
                 P
                 , 
                 
                 4606
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010111; B = 7'b1100001; // Expected: {'P': 8439}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010111; B = 7'b1100001; | Outputs: P=%b | Expected: P=%d",
                 2580,
                 
                 P
                 , 
                 
                 8439
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111110; B = 7'b0001000; // Expected: {'P': 1008}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111110; B = 7'b0001000; | Outputs: P=%b | Expected: P=%d",
                 2581,
                 
                 P
                 , 
                 
                 1008
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110010; B = 7'b0001100; // Expected: {'P': 1368}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110010; B = 7'b0001100; | Outputs: P=%b | Expected: P=%d",
                 2582,
                 
                 P
                 , 
                 
                 1368
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011101; B = 7'b0110011; // Expected: {'P': 1479}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011101; B = 7'b0110011; | Outputs: P=%b | Expected: P=%d",
                 2583,
                 
                 P
                 , 
                 
                 1479
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011111; B = 7'b1010101; // Expected: {'P': 8075}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011111; B = 7'b1010101; | Outputs: P=%b | Expected: P=%d",
                 2584,
                 
                 P
                 , 
                 
                 8075
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100011; B = 7'b1110011; // Expected: {'P': 4025}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100011; B = 7'b1110011; | Outputs: P=%b | Expected: P=%d",
                 2585,
                 
                 P
                 , 
                 
                 4025
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111100; B = 7'b1111101; // Expected: {'P': 7500}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111100; B = 7'b1111101; | Outputs: P=%b | Expected: P=%d",
                 2586,
                 
                 P
                 , 
                 
                 7500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001001; B = 7'b1100110; // Expected: {'P': 918}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001001; B = 7'b1100110; | Outputs: P=%b | Expected: P=%d",
                 2587,
                 
                 P
                 , 
                 
                 918
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100101; B = 7'b1011010; // Expected: {'P': 9090}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100101; B = 7'b1011010; | Outputs: P=%b | Expected: P=%d",
                 2588,
                 
                 P
                 , 
                 
                 9090
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010110; B = 7'b0110110; // Expected: {'P': 1188}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010110; B = 7'b0110110; | Outputs: P=%b | Expected: P=%d",
                 2589,
                 
                 P
                 , 
                 
                 1188
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110000; B = 7'b1011000; // Expected: {'P': 9856}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110000; B = 7'b1011000; | Outputs: P=%b | Expected: P=%d",
                 2590,
                 
                 P
                 , 
                 
                 9856
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111001; B = 7'b0110001; // Expected: {'P': 5929}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111001; B = 7'b0110001; | Outputs: P=%b | Expected: P=%d",
                 2591,
                 
                 P
                 , 
                 
                 5929
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000111; B = 7'b1010110; // Expected: {'P': 6106}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000111; B = 7'b1010110; | Outputs: P=%b | Expected: P=%d",
                 2592,
                 
                 P
                 , 
                 
                 6106
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000100; B = 7'b0111011; // Expected: {'P': 236}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000100; B = 7'b0111011; | Outputs: P=%b | Expected: P=%d",
                 2593,
                 
                 P
                 , 
                 
                 236
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000110; B = 7'b1010111; // Expected: {'P': 522}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000110; B = 7'b1010111; | Outputs: P=%b | Expected: P=%d",
                 2594,
                 
                 P
                 , 
                 
                 522
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000101; B = 7'b0000001; // Expected: {'P': 69}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000101; B = 7'b0000001; | Outputs: P=%b | Expected: P=%d",
                 2595,
                 
                 P
                 , 
                 
                 69
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101001; B = 7'b1111001; // Expected: {'P': 4961}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101001; B = 7'b1111001; | Outputs: P=%b | Expected: P=%d",
                 2596,
                 
                 P
                 , 
                 
                 4961
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001100; B = 7'b0010111; // Expected: {'P': 276}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001100; B = 7'b0010111; | Outputs: P=%b | Expected: P=%d",
                 2597,
                 
                 P
                 , 
                 
                 276
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000101; B = 7'b1111001; // Expected: {'P': 8349}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000101; B = 7'b1111001; | Outputs: P=%b | Expected: P=%d",
                 2598,
                 
                 P
                 , 
                 
                 8349
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000011; B = 7'b0100001; // Expected: {'P': 2211}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000011; B = 7'b0100001; | Outputs: P=%b | Expected: P=%d",
                 2599,
                 
                 P
                 , 
                 
                 2211
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111110; B = 7'b0001100; // Expected: {'P': 744}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111110; B = 7'b0001100; | Outputs: P=%b | Expected: P=%d",
                 2600,
                 
                 P
                 , 
                 
                 744
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000010; B = 7'b1010100; // Expected: {'P': 168}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000010; B = 7'b1010100; | Outputs: P=%b | Expected: P=%d",
                 2601,
                 
                 P
                 , 
                 
                 168
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100111; B = 7'b1111111; // Expected: {'P': 4953}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100111; B = 7'b1111111; | Outputs: P=%b | Expected: P=%d",
                 2602,
                 
                 P
                 , 
                 
                 4953
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001101; B = 7'b1001111; // Expected: {'P': 6083}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001101; B = 7'b1001111; | Outputs: P=%b | Expected: P=%d",
                 2603,
                 
                 P
                 , 
                 
                 6083
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100101; B = 7'b1110100; // Expected: {'P': 4292}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100101; B = 7'b1110100; | Outputs: P=%b | Expected: P=%d",
                 2604,
                 
                 P
                 , 
                 
                 4292
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001110; B = 7'b1011000; // Expected: {'P': 1232}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001110; B = 7'b1011000; | Outputs: P=%b | Expected: P=%d",
                 2605,
                 
                 P
                 , 
                 
                 1232
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011110; B = 7'b0001001; // Expected: {'P': 846}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011110; B = 7'b0001001; | Outputs: P=%b | Expected: P=%d",
                 2606,
                 
                 P
                 , 
                 
                 846
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111011; B = 7'b1001011; // Expected: {'P': 4425}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111011; B = 7'b1001011; | Outputs: P=%b | Expected: P=%d",
                 2607,
                 
                 P
                 , 
                 
                 4425
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100100; B = 7'b1110100; // Expected: {'P': 11600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100100; B = 7'b1110100; | Outputs: P=%b | Expected: P=%d",
                 2608,
                 
                 P
                 , 
                 
                 11600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001100; B = 7'b0101101; // Expected: {'P': 540}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001100; B = 7'b0101101; | Outputs: P=%b | Expected: P=%d",
                 2609,
                 
                 P
                 , 
                 
                 540
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010000; B = 7'b0010100; // Expected: {'P': 1600}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010000; B = 7'b0010100; | Outputs: P=%b | Expected: P=%d",
                 2610,
                 
                 P
                 , 
                 
                 1600
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011011; B = 7'b1100001; // Expected: {'P': 8827}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011011; B = 7'b1100001; | Outputs: P=%b | Expected: P=%d",
                 2611,
                 
                 P
                 , 
                 
                 8827
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011111; B = 7'b0001101; // Expected: {'P': 403}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011111; B = 7'b0001101; | Outputs: P=%b | Expected: P=%d",
                 2612,
                 
                 P
                 , 
                 
                 403
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000011; B = 7'b1000110; // Expected: {'P': 4690}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000011; B = 7'b1000110; | Outputs: P=%b | Expected: P=%d",
                 2613,
                 
                 P
                 , 
                 
                 4690
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010111; B = 7'b1011010; // Expected: {'P': 7830}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010111; B = 7'b1011010; | Outputs: P=%b | Expected: P=%d",
                 2614,
                 
                 P
                 , 
                 
                 7830
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100101; B = 7'b0001101; // Expected: {'P': 481}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100101; B = 7'b0001101; | Outputs: P=%b | Expected: P=%d",
                 2615,
                 
                 P
                 , 
                 
                 481
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110101; B = 7'b1100011; // Expected: {'P': 11583}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110101; B = 7'b1100011; | Outputs: P=%b | Expected: P=%d",
                 2616,
                 
                 P
                 , 
                 
                 11583
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111101; B = 7'b0000110; // Expected: {'P': 750}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111101; B = 7'b0000110; | Outputs: P=%b | Expected: P=%d",
                 2617,
                 
                 P
                 , 
                 
                 750
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000001; B = 7'b0011001; // Expected: {'P': 25}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000001; B = 7'b0011001; | Outputs: P=%b | Expected: P=%d",
                 2618,
                 
                 P
                 , 
                 
                 25
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110011; B = 7'b1101000; // Expected: {'P': 5304}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110011; B = 7'b1101000; | Outputs: P=%b | Expected: P=%d",
                 2619,
                 
                 P
                 , 
                 
                 5304
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000011; B = 7'b0101101; // Expected: {'P': 135}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000011; B = 7'b0101101; | Outputs: P=%b | Expected: P=%d",
                 2620,
                 
                 P
                 , 
                 
                 135
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111001; B = 7'b0100010; // Expected: {'P': 1938}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111001; B = 7'b0100010; | Outputs: P=%b | Expected: P=%d",
                 2621,
                 
                 P
                 , 
                 
                 1938
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100011; B = 7'b1101000; // Expected: {'P': 10296}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100011; B = 7'b1101000; | Outputs: P=%b | Expected: P=%d",
                 2622,
                 
                 P
                 , 
                 
                 10296
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011110; B = 7'b0100010; // Expected: {'P': 1020}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011110; B = 7'b0100010; | Outputs: P=%b | Expected: P=%d",
                 2623,
                 
                 P
                 , 
                 
                 1020
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101110; B = 7'b1011001; // Expected: {'P': 4094}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101110; B = 7'b1011001; | Outputs: P=%b | Expected: P=%d",
                 2624,
                 
                 P
                 , 
                 
                 4094
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110011; B = 7'b1001100; // Expected: {'P': 8740}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110011; B = 7'b1001100; | Outputs: P=%b | Expected: P=%d",
                 2625,
                 
                 P
                 , 
                 
                 8740
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000101; B = 7'b1101000; // Expected: {'P': 520}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000101; B = 7'b1101000; | Outputs: P=%b | Expected: P=%d",
                 2626,
                 
                 P
                 , 
                 
                 520
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001101; B = 7'b0110110; // Expected: {'P': 702}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001101; B = 7'b0110110; | Outputs: P=%b | Expected: P=%d",
                 2627,
                 
                 P
                 , 
                 
                 702
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011001; B = 7'b1010001; // Expected: {'P': 7209}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011001; B = 7'b1010001; | Outputs: P=%b | Expected: P=%d",
                 2628,
                 
                 P
                 , 
                 
                 7209
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001011; B = 7'b0010100; // Expected: {'P': 1500}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001011; B = 7'b0010100; | Outputs: P=%b | Expected: P=%d",
                 2629,
                 
                 P
                 , 
                 
                 1500
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011100; B = 7'b0110110; // Expected: {'P': 4968}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011100; B = 7'b0110110; | Outputs: P=%b | Expected: P=%d",
                 2630,
                 
                 P
                 , 
                 
                 4968
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010011; B = 7'b0101101; // Expected: {'P': 3735}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010011; B = 7'b0101101; | Outputs: P=%b | Expected: P=%d",
                 2631,
                 
                 P
                 , 
                 
                 3735
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110110; B = 7'b1011001; // Expected: {'P': 10502}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110110; B = 7'b1011001; | Outputs: P=%b | Expected: P=%d",
                 2632,
                 
                 P
                 , 
                 
                 10502
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1111001; B = 7'b1100111; // Expected: {'P': 12463}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1111001; B = 7'b1100111; | Outputs: P=%b | Expected: P=%d",
                 2633,
                 
                 P
                 , 
                 
                 12463
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011001; B = 7'b0111101; // Expected: {'P': 5429}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011001; B = 7'b0111101; | Outputs: P=%b | Expected: P=%d",
                 2634,
                 
                 P
                 , 
                 
                 5429
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011000; B = 7'b1000100; // Expected: {'P': 1632}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011000; B = 7'b1000100; | Outputs: P=%b | Expected: P=%d",
                 2635,
                 
                 P
                 , 
                 
                 1632
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111101; B = 7'b1111010; // Expected: {'P': 7442}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111101; B = 7'b1111010; | Outputs: P=%b | Expected: P=%d",
                 2636,
                 
                 P
                 , 
                 
                 7442
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000110; B = 7'b0011110; // Expected: {'P': 180}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000110; B = 7'b0011110; | Outputs: P=%b | Expected: P=%d",
                 2637,
                 
                 P
                 , 
                 
                 180
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1110101; B = 7'b1010100; // Expected: {'P': 9828}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1110101; B = 7'b1010100; | Outputs: P=%b | Expected: P=%d",
                 2638,
                 
                 P
                 , 
                 
                 9828
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110001; B = 7'b1001000; // Expected: {'P': 3528}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110001; B = 7'b1001000; | Outputs: P=%b | Expected: P=%d",
                 2639,
                 
                 P
                 , 
                 
                 3528
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110000; B = 7'b0011111; // Expected: {'P': 1488}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110000; B = 7'b0011111; | Outputs: P=%b | Expected: P=%d",
                 2640,
                 
                 P
                 , 
                 
                 1488
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111010; B = 7'b1001101; // Expected: {'P': 4466}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111010; B = 7'b1001101; | Outputs: P=%b | Expected: P=%d",
                 2641,
                 
                 P
                 , 
                 
                 4466
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001001; B = 7'b0011001; // Expected: {'P': 225}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001001; B = 7'b0011001; | Outputs: P=%b | Expected: P=%d",
                 2642,
                 
                 P
                 , 
                 
                 225
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0011000; B = 7'b1101000; // Expected: {'P': 2496}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0011000; B = 7'b1101000; | Outputs: P=%b | Expected: P=%d",
                 2643,
                 
                 P
                 , 
                 
                 2496
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0001111; B = 7'b0101010; // Expected: {'P': 630}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0001111; B = 7'b0101010; | Outputs: P=%b | Expected: P=%d",
                 2644,
                 
                 P
                 , 
                 
                 630
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111001; B = 7'b1010101; // Expected: {'P': 4845}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111001; B = 7'b1010101; | Outputs: P=%b | Expected: P=%d",
                 2645,
                 
                 P
                 , 
                 
                 4845
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001000; B = 7'b1011011; // Expected: {'P': 6552}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001000; B = 7'b1011011; | Outputs: P=%b | Expected: P=%d",
                 2646,
                 
                 P
                 , 
                 
                 6552
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1000100; B = 7'b0101001; // Expected: {'P': 2788}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1000100; B = 7'b0101001; | Outputs: P=%b | Expected: P=%d",
                 2647,
                 
                 P
                 , 
                 
                 2788
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0000000; B = 7'b1010010; // Expected: {'P': 0}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0000000; B = 7'b1010010; | Outputs: P=%b | Expected: P=%d",
                 2648,
                 
                 P
                 , 
                 
                 0
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101100; B = 7'b1000100; // Expected: {'P': 2992}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101100; B = 7'b1000100; | Outputs: P=%b | Expected: P=%d",
                 2649,
                 
                 P
                 , 
                 
                 2992
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0010000; B = 7'b0011001; // Expected: {'P': 400}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0010000; B = 7'b0011001; | Outputs: P=%b | Expected: P=%d",
                 2650,
                 
                 P
                 , 
                 
                 400
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1100101; B = 7'b0100001; // Expected: {'P': 3333}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1100101; B = 7'b0100001; | Outputs: P=%b | Expected: P=%d",
                 2651,
                 
                 P
                 , 
                 
                 3333
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011101; B = 7'b1101111; // Expected: {'P': 10323}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011101; B = 7'b1101111; | Outputs: P=%b | Expected: P=%d",
                 2652,
                 
                 P
                 , 
                 
                 10323
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1001010; B = 7'b0100001; // Expected: {'P': 2442}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1001010; B = 7'b0100001; | Outputs: P=%b | Expected: P=%d",
                 2653,
                 
                 P
                 , 
                 
                 2442
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0100110; B = 7'b1100010; // Expected: {'P': 3724}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0100110; B = 7'b1100010; | Outputs: P=%b | Expected: P=%d",
                 2654,
                 
                 P
                 , 
                 
                 3724
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1011111; B = 7'b1001110; // Expected: {'P': 7410}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1011111; B = 7'b1001110; | Outputs: P=%b | Expected: P=%d",
                 2655,
                 
                 P
                 , 
                 
                 7410
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0111101; B = 7'b1011100; // Expected: {'P': 5612}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0111101; B = 7'b1011100; | Outputs: P=%b | Expected: P=%d",
                 2656,
                 
                 P
                 , 
                 
                 5612
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b1010110; B = 7'b0111101; // Expected: {'P': 5246}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b1010110; B = 7'b0111101; | Outputs: P=%b | Expected: P=%d",
                 2657,
                 
                 P
                 , 
                 
                 5246
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0110010; B = 7'b1110101; // Expected: {'P': 5850}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0110010; B = 7'b1110101; | Outputs: P=%b | Expected: P=%d",
                 2658,
                 
                 P
                 , 
                 
                 5850
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        #10 A = 7'b0101000; B = 7'b0011110; // Expected: {'P': 1200}
        
        
        #10;
        
        
        $display("Test %0d: Inputs: A = 7'b0101000; B = 7'b0011110; | Outputs: P=%b | Expected: P=%d",
                 2659,
                 
                 P
                 , 
                 
                 1200
                 
        );
        $timeformat(-9, 1, " ns", 6);
        $display("Simulation time: %t", $time);
        
        $finish;
    end
  
endmodule